CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
130 100 1 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
110
9 2-In AND~
219 784 1661 0 1 22
0 0
0
0 0 608 270
5 74F08
-18 -24 17 -16
4 U22A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5130 0 0
2
42660.2 0
0
13 Logic Switch~
5 332 1289 0 10 11
0 104 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V31
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
391 0 0
2
5.89773e-315 5.32571e-315
0
13 Logic Switch~
5 365 1291 0 1 11
0 105
0
0 0 21360 90
2 0V
11 0 25 8
3 V30
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -2 0
1 V
3124 0 0
2
5.89773e-315 5.30499e-315
0
13 Logic Switch~
5 396 1291 0 1 11
0 106
0
0 0 21360 90
2 0V
11 0 25 8
3 V29
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -2 0
1 V
3421 0 0
2
5.89773e-315 5.26354e-315
0
13 Logic Switch~
5 428 1292 0 1 11
0 107
0
0 0 21360 90
2 0V
11 0 25 8
3 V28
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -2 0
1 V
8157 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1701 375 0 1 11
0 36
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V41
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1707 634 0 1 11
0 45
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V40
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1742 556 0 1 11
0 49
0
0 0 21360 90
2 0V
11 0 25 8
3 V39
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.89773e-315 5.32571e-315
0
13 Logic Switch~
5 1775 558 0 1 11
0 48
0
0 0 21360 90
2 0V
11 0 25 8
3 V38
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.89773e-315 5.30499e-315
0
13 Logic Switch~
5 1806 558 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V37
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.89773e-315 5.26354e-315
0
13 Logic Switch~
5 1838 559 0 1 11
0 46
0
0 0 21360 90
2 0V
11 0 25 8
3 V36
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 101 110 0 1 11
0 54
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V27
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 102 295 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 105 564 0 10 11
0 63 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V25
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 380 501 0 10 11
0 70 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V20
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.89773e-315 5.32571e-315
0
13 Logic Switch~
5 348 500 0 1 11
0 71
0
0 0 21360 90
2 0V
11 0 25 8
3 V22
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3670 0 0
2
5.89773e-315 5.30499e-315
0
13 Logic Switch~
5 317 500 0 10 11
0 72 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V23
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.89773e-315 5.26354e-315
0
13 Logic Switch~
5 284 498 0 10 11
0 73 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V24
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 103 359 0 10 11
0 69 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 101 158 0 10 11
0 74 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3108 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 100 68 0 1 11
0 76
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4299 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 101 1238 0 1 11
0 86
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9672 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 104 1059 0 1 11
0 91
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7876 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1708 1033 0 1 11
0 96
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V14
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1709 802 0 1 11
0 81
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V13
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9172 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1536 965 0 1 11
0 100
0
0 0 21360 90
2 0V
11 0 25 8
3 V12
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
5.89773e-315 5.32571e-315
0
13 Logic Switch~
5 1569 967 0 1 11
0 99
0
0 0 21360 90
2 0V
11 0 25 8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3820 0 0
2
5.89773e-315 5.30499e-315
0
13 Logic Switch~
5 1600 967 0 1 11
0 98
0
0 0 21360 90
2 0V
11 0 25 8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
5.89773e-315 5.26354e-315
0
13 Logic Switch~
5 1632 968 0 1 11
0 97
0
0 0 21360 90
2 0V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1385 966 0 10 11
0 85 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1353 965 0 1 11
0 84
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1322 965 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3951 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1289 963 0 10 11
0 82 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1708 762 0 1 11
0 101
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1700 325 0 1 11
0 102
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9265 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 1696 141 0 1 11
0 103
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9442 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 100 31 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
5.89773e-315 0
0
2 +V
167 675 1372 0 1 3
0 4
0
0 0 54256 180
3 10V
6 -2 27 6
3 V32
6 -12 27 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9968 0 0
2
42660.2 0
0
9 3-In NOR~
219 711 1261 0 4 22
0 7 6 5 8
0
0 0 624 180
5 74F27
-18 -24 17 -16
4 U21A
-11 -2 17 6
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
9281 0 0
2
42660.2 0
0
14 Logic Display~
6 1552 1300 0 1 2
10 5
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L33
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
42660.2 3
0
14 Logic Display~
6 1552 1325 0 1 2
10 6
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L32
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
42660.2 2
0
14 Logic Display~
6 1552 1351 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L31
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
42660.2 1
0
14 Logic Display~
6 1552 1274 0 1 2
10 9
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L30
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
42660.2 0
0
7 74LS164
127 716 1324 0 12 25
0 8 8 3 4 108 109 110 111 9
5 6 7
0
0 0 4848 0
6 74F164
-21 -51 21 -43
3 U20
-14 4 7 12
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 512 0 0 0 0
1 U
6435 0 0
2
42660.2 0
0
14 Logic Display~
6 1550 1405 0 1 2
10 18
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L21
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.89773e-315 5.38788e-315
0
14 Logic Display~
6 1550 1482 0 1 2
10 15
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L23
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
5.89773e-315 5.37752e-315
0
14 Logic Display~
6 1550 1456 0 1 2
10 16
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L24
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.89773e-315 5.36716e-315
0
14 Logic Display~
6 1549 1558 0 1 2
10 12
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L25
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.89773e-315 5.3568e-315
0
14 Logic Display~
6 1550 1584 0 1 2
10 11
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L26
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.89773e-315 5.34643e-315
0
14 Logic Display~
6 1549 1533 0 1 2
10 13
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L27
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.89773e-315 5.32571e-315
0
14 Logic Display~
6 1549 1507 0 1 2
10 14
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L28
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.89773e-315 5.30499e-315
0
14 Logic Display~
6 1550 1608 0 1 2
10 10
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L29
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.89773e-315 5.26354e-315
0
14 Logic Display~
6 1550 1431 0 1 2
10 17
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.89773e-315 0
0
9 Inverter~
13 662 1610 0 2 22
0 19 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
34 0 0
2
5.89773e-315 5.26354e-315
0
9 Inverter~
13 662 1509 0 2 22
0 23 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
6357 0 0
2
5.89773e-315 5.32571e-315
0
9 Inverter~
13 662 1535 0 2 22
0 22 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
319 0 0
2
5.89773e-315 5.30499e-315
0
9 Inverter~
13 662 1586 0 2 22
0 20 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3976 0 0
2
5.89773e-315 5.26354e-315
0
9 Inverter~
13 662 1560 0 2 22
0 21 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
7634 0 0
2
5.89773e-315 0
0
9 Inverter~
13 663 1458 0 2 22
0 25 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
523 0 0
2
5.89773e-315 5.26354e-315
0
9 Inverter~
13 663 1484 0 2 22
0 24 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
6748 0 0
2
5.89773e-315 0
0
9 Inverter~
13 663 1433 0 2 22
0 26 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
6901 0 0
2
5.89773e-315 0
0
9 Inverter~
13 663 1407 0 2 22
0 27 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
842 0 0
2
5.89773e-315 0
0
7 Ground~
168 586 1270 0 1 3
0 2
0
0 0 53360 90
0
5 GND10
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3277 0 0
2
5.89773e-315 0
0
7 74LS154
95 551 1316 0 22 45
0 2 2 28 29 30 31 112 113 114
115 116 117 118 19 20 21 22 23 24
25 26 27
0
0 0 4848 270
6 74F154
-21 -87 21 -79
3 U17
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
4212 0 0
2
5.89773e-315 0
0
9 4-In NOR~
219 1422 275 0 5 22
0 35 34 33 32 119
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 1 1 0
1 U
4720 0 0
2
5.89773e-315 0
0
7 74LS126
116 1089 430 0 12 25
0 36 37 36 38 36 39 36 40 41
42 43 44
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
3 U15
-10 -52 11 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
5551 0 0
2
5.89773e-315 0
0
7 Ground~
168 1108 510 0 1 3
0 2
0
0 0 53360 270
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6986 0 0
2
5.89773e-315 0
0
7 74LS181
132 1190 471 0 22 45
0 49 48 47 46 32 33 34 35 53
52 51 50 45 2 120 121 122 123 37
38 39 40
0
0 0 4848 180
7 74LS181
-24 -69 25 -61
3 U14
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
8745 0 0
2
5.89773e-315 0
0
6 PROM32
80 777 600 0 14 29
0 63 2 62 61 60 59 55 56 57
58 41 42 43 44
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9592 0 0
2
5.89773e-315 0
0
BBFFIIAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 Ground~
168 389 599 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8748 0 0
2
5.89773e-315 0
0
7 74LS173
129 771 440 0 14 29
0 2 68 68 3 44 43 42 41 2
2 64 65 66 67
0
0 0 4848 270
6 74F173
-21 -51 21 -43
3 U12
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
5.89773e-315 5.26354e-315
0
7 Ground~
168 869 405 0 1 3
0 2
0
0 0 53360 90
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
631 0 0
2
5.89773e-315 0
0
7 Ground~
168 546 479 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9466 0 0
2
5.89773e-315 0
0
7 74LS257
147 614 517 0 14 29
0 69 64 70 65 71 66 72 67 73
2 59 60 61 62
0
0 0 4848 270
6 74F257
-21 -60 21 -52
3 U11
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3266 0 0
2
5.89773e-315 0
0
7 Ground~
168 475 168 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7693 0 0
2
5.89773e-315 0
0
2 +V
167 598 114 0 1 3
0 75
0
0 0 54256 0
2 5V
-8 -22 6 -14
3 V17
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3723 0 0
2
5.89773e-315 0
0
7 74LS193
137 663 168 0 14 29
0 54 75 74 2 41 42 43 44 124
125 80 79 78 77
0
0 0 4848 0
6 74F193
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3440 0 0
2
5.89773e-315 0
0
7 74LS126
116 826 169 0 12 25
0 76 80 76 79 76 78 76 77 41
42 43 44
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
6263 0 0
2
5.89773e-315 0
0
7 74LS126
116 845 1176 0 12 25
0 86 87 86 88 86 89 86 90 44
43 42 41
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U8
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
4900 0 0
2
5.89773e-315 0
0
7 Ground~
168 743 1174 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8783 0 0
2
5.89773e-315 0
0
7 74LS173
129 671 1128 0 14 29
0 2 91 91 3 44 43 42 41 2
2 87 88 89 90
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U7
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3221 0 0
2
5.89773e-315 0
0
7 74LS173
129 542 1127 0 14 29
0 2 91 91 3 58 57 56 55 2
2 28 29 30 31
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U6
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3215 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 1390 1160 0 1 2
10 95
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
5.89773e-315 5.32571e-315
0
14 Logic Display~
6 1370 1160 0 1 2
10 94
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7121 0 0
2
5.89773e-315 5.30499e-315
0
14 Logic Display~
6 1350 1160 0 1 2
10 93
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
5.89773e-315 5.26354e-315
0
14 Logic Display~
6 1331 1160 0 1 2
10 92
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.89773e-315 0
0
7 Ground~
168 1253 1131 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7804 0 0
2
5.89773e-315 0
0
7 74LS173
129 1158 1090 0 14 29
0 2 96 96 3 41 42 43 44 2
2 92 93 94 95
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U5
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
5523 0 0
2
5.89773e-315 0
0
7 Ground~
168 1400 746 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3330 0 0
2
5.89773e-315 0
0
7 74LS126
116 1090 852 0 12 25
0 81 82 81 83 81 84 81 85 41
42 43 44
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3465 0 0
2
5.89773e-315 0
0
7 74LS257
147 1323 708 0 14 29
0 101 82 100 83 99 84 98 85 97
2 53 52 51 50
0
0 0 4848 90
6 74F257
-21 -60 21 -52
2 U3
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8396 0 0
2
5.89773e-315 0
0
7 74LS126
116 1091 294 0 12 25
0 102 32 102 33 102 34 102 35 41
42 43 44
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3685 0 0
2
5.89773e-315 0
0
7 Ground~
168 1254 242 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7849 0 0
2
5.89773e-315 0
0
7 74LS173
129 1159 200 0 14 29
0 2 103 103 3 41 42 43 44 2
2 32 33 34 35
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U1
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6343 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 916 1239 0 1 2
10 55
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L16
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
42660.1 0
0
14 Logic Display~
6 935 1239 0 1 2
10 56
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L15
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
42660.1 1
0
14 Logic Display~
6 955 1239 0 1 2
10 57
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L14
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
42660.1 2
0
14 Logic Display~
6 975 1239 0 1 2
10 58
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L13
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
42660.1 3
0
14 Logic Display~
6 1053 1239 0 1 2
10 44
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L12
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
42660.1 4
0
14 Logic Display~
6 1033 1239 0 1 2
10 43
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L11
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
42660.1 5
0
14 Logic Display~
6 1013 1239 0 1 2
10 42
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L10
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
42660.1 6
0
14 Logic Display~
6 994 1239 0 1 2
10 41
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
42660.1 7
0
14 Logic Display~
6 994 94 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7978 0 0
2
42660.1 8
0
14 Logic Display~
6 1013 94 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3142 0 0
2
42660.1 9
0
14 Logic Display~
6 1033 94 0 1 2
10 43
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
42660.1 10
0
14 Logic Display~
6 1053 94 0 1 2
10 44
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
659 0 0
2
42660.1 11
0
14 Logic Display~
6 975 94 0 1 2
10 58
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
42660.1 12
0
14 Logic Display~
6 955 94 0 1 2
10 57
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6792 0 0
2
42660.1 13
0
14 Logic Display~
6 935 94 0 1 2
10 56
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
42660.1 14
0
14 Logic Display~
6 916 94 0 1 2
10 55
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6316 0 0
2
42660.1 15
0
220
1 5 0 0 0 0 0 1 65 0 0 5
791 1639
791 1260
1486 1260
1486 275
1461 275
2 0 0 0 0 0 0 1 0 0 15 2
773 1639
773 1588
3 0 3 0 0 12288 0 44 0 0 163 5
684 1324
659 1324
659 1225
167 1225
167 1020
1 4 4 0 0 8320 0 38 44 0 0 3
675 1357
678 1357
678 1342
3 0 5 0 0 8192 0 39 0 0 11 3
736 1252
779 1252
779 1304
2 0 6 0 0 8192 0 39 0 0 12 3
735 1261
774 1261
774 1329
1 0 7 0 0 8192 0 39 0 0 13 3
736 1270
770 1270
770 1355
2 0 8 0 0 4096 0 44 0 0 9 3
684 1306
669 1306
669 1297
1 4 8 0 0 8320 0 44 39 0 0 4
684 1297
669 1297
669 1261
684 1261
9 1 9 0 0 12416 0 44 43 0 0 4
748 1333
766 1333
766 1278
1536 1278
10 1 5 0 0 12416 0 44 40 0 0 4
748 1342
759 1342
759 1304
1536 1304
1 11 6 0 0 4224 0 41 44 0 0 4
1536 1329
754 1329
754 1351
748 1351
1 12 7 0 0 4224 0 42 44 0 0 4
1536 1355
754 1355
754 1360
748 1360
2 1 10 0 0 8320 0 54 52 0 0 3
683 1610
683 1612
1534 1612
2 1 11 0 0 8320 0 57 49 0 0 3
683 1586
683 1588
1534 1588
2 1 12 0 0 8320 0 58 48 0 0 3
683 1560
683 1562
1533 1562
2 1 13 0 0 8320 0 56 50 0 0 3
683 1535
683 1537
1533 1537
2 1 14 0 0 8320 0 55 51 0 0 3
683 1509
683 1511
1533 1511
2 1 15 0 0 8320 0 60 46 0 0 3
684 1484
684 1486
1534 1486
2 1 16 0 0 8320 0 59 47 0 0 3
684 1458
684 1460
1534 1460
2 1 17 0 0 8320 0 61 53 0 0 3
684 1433
684 1435
1534 1435
2 1 18 0 0 8320 0 62 45 0 0 3
684 1407
684 1409
1534 1409
0 2 10 0 0 0 0 0 54 0 0 4
684 1610
682 1610
682 1610
683 1610
14 1 19 0 0 4224 0 64 54 0 0 3
553 1356
553 1610
647 1610
15 1 20 0 0 4224 0 64 57 0 0 3
544 1356
544 1586
647 1586
1 16 21 0 0 8320 0 58 64 0 0 3
647 1560
535 1560
535 1356
17 1 22 0 0 4224 0 64 56 0 0 3
526 1356
526 1535
647 1535
18 1 23 0 0 4224 0 64 55 0 0 3
517 1356
517 1509
647 1509
19 1 24 0 0 8320 0 64 60 0 0 3
508 1356
508 1484
648 1484
20 1 25 0 0 8320 0 64 59 0 0 3
499 1356
499 1458
648 1458
21 1 26 0 0 8320 0 64 61 0 0 3
490 1356
490 1433
648 1433
22 1 27 0 0 8320 0 64 62 0 0 3
481 1356
481 1407
648 1407
1 0 2 0 0 4096 0 64 0 0 34 2
571 1280
571 1271
1 2 2 0 0 4096 0 63 64 0 0 3
579 1271
562 1271
562 1280
11 3 28 0 0 4224 0 82 64 0 0 2
535 1161
535 1286
12 4 29 0 0 4224 0 82 64 0 0 2
526 1161
526 1286
13 5 30 0 0 4224 0 82 64 0 0 2
517 1161
517 1286
6 14 31 0 0 4224 0 64 82 0 0 2
508 1286
508 1161
0 4 32 0 0 4096 0 0 65 46 0 4
1233 316
1356 316
1356 289
1405 289
0 3 33 0 0 4096 0 0 65 45 0 4
1245 299
1343 299
1343 280
1405 280
0 2 34 0 0 4096 0 0 65 44 0 4
1255 282
1334 282
1334 271
1405 271
0 1 35 0 0 4096 0 0 65 43 0 2
1265 262
1405 262
8 8 35 0 0 8320 0 68 92 0 0 4
1228 457
1265 457
1265 262
1123 262
7 0 34 0 0 8320 0 68 0 0 201 4
1228 466
1255 466
1255 280
1134 280
6 0 33 0 0 8320 0 68 0 0 200 4
1228 475
1245 475
1245 298
1143 298
0 5 32 0 0 8320 0 0 68 199 0 4
1152 316
1236 316
1236 484
1228 484
7 0 36 0 0 4096 0 66 0 0 50 2
1121 407
1128 407
5 0 36 0 0 0 0 66 0 0 50 2
1121 425
1128 425
3 0 36 0 0 0 0 66 0 0 50 2
1121 443
1128 443
1 1 36 0 0 4224 0 6 66 0 0 4
1687 375
1128 375
1128 461
1121 461
2 19 37 0 0 4224 0 66 68 0 0 3
1121 452
1152 452
1152 448
4 20 38 0 0 4224 0 66 68 0 0 4
1121 434
1147 434
1147 439
1152 439
6 21 39 0 0 4224 0 66 68 0 0 4
1121 416
1142 416
1142 430
1152 430
22 8 40 0 0 12416 0 68 66 0 0 4
1152 421
1146 421
1146 398
1121 398
9 0 41 0 0 4096 0 66 0 0 216 2
1057 452
994 452
10 0 42 0 0 4096 0 66 0 0 215 2
1057 434
1013 434
11 0 43 0 0 4096 0 66 0 0 214 2
1057 416
1033 416
12 0 44 0 0 4096 0 66 0 0 213 2
1057 398
1053 398
14 1 2 0 0 4096 0 68 67 0 0 2
1158 511
1115 511
13 1 45 0 0 12416 0 68 7 0 0 4
1158 520
1146 520
1146 634
1693 634
4 1 46 0 0 4224 0 68 11 0 0 3
1222 493
1839 493
1839 546
3 1 47 0 0 4224 0 68 10 0 0 3
1222 502
1807 502
1807 545
2 1 48 0 0 4224 0 68 9 0 0 3
1222 511
1776 511
1776 545
1 1 49 0 0 4224 0 68 8 0 0 3
1222 520
1743 520
1743 543
12 14 50 0 0 8320 0 68 91 0 0 3
1228 421
1354 421
1354 675
11 13 51 0 0 8320 0 68 91 0 0 3
1228 430
1336 430
1336 675
10 12 52 0 0 8320 0 68 91 0 0 3
1228 439
1318 439
1318 675
9 11 53 0 0 8320 0 68 91 0 0 3
1228 448
1300 448
1300 675
1 1 54 0 0 4224 0 12 77 0 0 4
113 110
385 110
385 141
631 141
8 0 55 0 0 8192 0 82 0 0 220 3
508 1097
508 935
916 935
0 7 56 0 0 4096 0 0 82 219 0 3
935 946
517 946
517 1097
6 0 57 0 0 8192 0 82 0 0 218 3
526 1097
526 961
955 961
5 0 58 0 0 8192 0 82 0 0 217 3
535 1097
535 975
975 975
11 6 59 0 0 8320 0 74 69 0 0 3
631 554
631 636
745 636
5 12 60 0 0 4224 0 69 74 0 0 3
745 627
613 627
613 554
13 4 61 0 0 8320 0 74 69 0 0 3
595 554
595 618
745 618
14 3 62 0 0 8320 0 74 69 0 0 3
577 554
577 609
745 609
14 0 44 0 0 4096 0 69 0 0 213 2
809 636
1053 636
13 0 43 0 0 4096 0 69 0 0 214 2
809 627
1033 627
12 0 42 0 0 4096 0 69 0 0 215 2
809 618
1013 618
11 0 41 0 0 4096 0 69 0 0 216 2
809 609
994 609
10 0 58 0 0 0 0 69 0 0 217 2
809 600
975 600
9 0 57 0 0 0 0 69 0 0 218 2
809 591
955 591
8 0 56 0 0 0 0 69 0 0 219 2
809 582
935 582
7 0 55 0 0 0 0 69 0 0 220 2
809 573
916 573
1 2 2 0 0 4224 0 70 69 0 0 2
396 600
745 600
1 1 63 0 0 4224 0 14 69 0 0 2
117 564
739 564
2 11 64 0 0 8320 0 74 71 0 0 4
640 490
640 483
764 483
764 474
12 4 65 0 0 8320 0 71 74 0 0 4
755 474
755 480
622 480
622 490
6 13 66 0 0 8320 0 74 71 0 0 4
604 490
604 477
746 477
746 474
14 8 67 0 0 4224 0 71 74 0 0 3
737 474
586 474
586 490
4 0 3 0 0 8192 0 71 0 0 163 3
773 410
773 275
167 275
5 0 44 0 0 8192 0 71 0 0 213 3
764 410
764 363
1053 363
6 0 43 0 0 8192 0 71 0 0 214 3
755 410
755 353
1033 353
7 0 42 0 0 8192 0 71 0 0 215 3
746 410
746 342
1013 342
8 0 41 0 0 8192 0 71 0 0 216 3
737 410
737 330
994 330
3 0 68 0 0 4096 0 71 0 0 98 3
782 404
782 395
791 395
1 2 68 0 0 4224 0 13 71 0 0 3
114 295
791 295
791 404
9 0 2 0 0 0 0 71 0 0 100 2
800 480
800 490
10 0 2 0 0 0 0 71 0 0 101 4
791 480
791 490
851 490
851 406
1 1 2 0 0 0 0 71 72 0 0 3
800 410
800 406
862 406
1 10 2 0 0 0 0 73 74 0 0 3
553 480
568 480
568 484
1 1 69 0 0 8320 0 74 19 0 0 3
649 490
649 359
115 359
1 3 70 0 0 8320 0 15 74 0 0 4
381 488
381 412
631 412
631 490
1 5 71 0 0 8320 0 16 74 0 0 4
349 487
349 397
613 397
613 490
1 7 72 0 0 8320 0 17 74 0 0 4
318 487
318 383
595 383
595 490
1 9 73 0 0 8320 0 18 74 0 0 4
285 485
285 370
577 370
577 490
9 0 41 0 0 0 0 78 0 0 216 2
858 151
994 151
10 0 42 0 0 0 0 78 0 0 215 2
858 169
1013 169
11 0 43 0 0 0 0 78 0 0 214 2
858 187
1033 187
12 0 44 0 0 0 0 78 0 0 213 2
858 205
1053 205
1 4 2 0 0 0 0 75 77 0 0 3
482 169
482 168
631 168
3 1 74 0 0 8320 0 77 20 0 0 3
625 159
625 158
113 158
2 1 75 0 0 4224 0 77 76 0 0 3
631 150
598 150
598 123
0 5 41 0 0 4096 0 0 77 216 0 4
994 248
593 248
593 177
631 177
0 6 42 0 0 4096 0 0 77 215 0 4
1013 240
602 240
602 186
631 186
0 7 43 0 0 4096 0 0 77 214 0 4
1033 231
611 231
611 195
631 195
0 8 44 0 0 4096 0 0 77 213 0 4
1053 222
620 222
620 204
631 204
1 0 76 0 0 4096 0 78 0 0 122 2
794 142
780 142
3 0 76 0 0 0 0 78 0 0 122 2
794 160
780 160
5 0 76 0 0 0 0 78 0 0 122 2
794 178
780 178
1 7 76 0 0 4224 0 21 78 0 0 4
112 68
780 68
780 196
794 196
8 14 77 0 0 8320 0 78 77 0 0 3
794 205
794 204
695 204
6 13 78 0 0 12416 0 78 77 0 0 4
794 187
748 187
748 195
695 195
4 12 79 0 0 4224 0 78 77 0 0 4
794 169
740 169
740 186
695 186
11 2 80 0 0 12416 0 77 78 0 0 4
695 177
731 177
731 151
794 151
7 0 81 0 0 4096 0 90 0 0 130 2
1122 829
1148 829
5 0 81 0 0 0 0 90 0 0 130 2
1122 847
1148 847
3 0 81 0 0 0 0 90 0 0 130 2
1122 865
1148 865
1 1 81 0 0 4224 0 25 90 0 0 4
1695 802
1148 802
1148 883
1122 883
2 0 82 0 0 4096 0 90 0 0 189 2
1122 874
1290 874
4 0 83 0 0 4096 0 90 0 0 188 2
1122 856
1309 856
6 0 84 0 0 4224 0 90 0 0 187 2
1122 838
1327 838
8 0 85 0 0 4224 0 90 0 0 186 2
1122 820
1345 820
7 0 86 0 0 4096 0 79 0 0 138 2
813 1203
758 1203
5 0 86 0 0 0 0 79 0 0 138 3
813 1185
813 1171
758 1171
3 0 86 0 0 0 0 79 0 0 138 2
813 1167
758 1167
1 1 86 0 0 4224 0 22 79 0 0 4
113 1238
758 1238
758 1149
813 1149
11 2 87 0 0 8320 0 81 79 0 0 5
664 1162
664 1186
793 1186
793 1158
813 1158
12 0 41 0 0 0 0 79 0 0 216 2
877 1212
994 1212
11 0 42 0 0 0 0 79 0 0 215 2
877 1194
1013 1194
10 0 43 0 0 0 0 79 0 0 214 2
877 1176
1033 1176
9 0 44 0 0 0 0 79 0 0 213 2
877 1158
1053 1158
12 4 88 0 0 8320 0 81 79 0 0 5
655 1162
655 1190
807 1190
807 1176
813 1176
13 6 89 0 0 8320 0 81 79 0 0 3
646 1162
646 1194
813 1194
14 8 90 0 0 8320 0 81 79 0 0 3
637 1162
637 1212
813 1212
3 0 91 0 0 8192 0 81 0 0 148 3
682 1092
682 1075
562 1075
1 2 91 0 0 4224 0 23 82 0 0 3
116 1059
562 1059
562 1091
3 2 91 0 0 0 0 82 82 0 0 2
553 1091
562 1091
3 2 91 0 0 0 0 81 81 0 0 2
682 1092
691 1092
0 0 3 0 0 0 0 0 0 152 163 2
673 1087
673 1020
4 4 3 0 0 0 0 81 82 0 0 4
673 1098
673 1085
544 1085
544 1097
1 0 2 0 0 0 0 80 0 0 154 4
736 1175
737 1175
737 1175
736 1175
1 0 2 0 0 0 0 81 0 0 155 4
700 1098
736 1098
736 1175
699 1175
0 9 2 0 0 0 0 0 81 156 0 3
690 1175
700 1175
700 1168
0 10 2 0 0 0 0 0 81 158 0 3
604 1175
691 1175
691 1168
9 0 2 0 0 0 0 82 0 0 158 2
571 1167
571 1176
1 10 2 0 0 0 0 82 82 0 0 5
571 1097
604 1097
604 1176
562 1176
562 1167
5 0 44 0 0 0 0 81 0 0 213 3
664 1098
664 1068
1053 1068
6 0 43 0 0 0 0 81 0 0 214 3
655 1098
655 1063
1033 1063
7 0 42 0 0 0 0 81 0 0 215 3
646 1098
646 1057
1013 1057
8 0 41 0 0 0 0 81 0 0 216 3
637 1098
637 1051
994 1051
4 0 3 0 0 8192 0 88 0 0 208 4
1160 1060
1160 1020
167 1020
167 31
11 1 92 0 0 8320 0 88 86 0 0 4
1151 1124
1151 1217
1331 1217
1331 1178
12 1 93 0 0 8320 0 88 85 0 0 4
1142 1124
1142 1210
1350 1210
1350 1178
13 1 94 0 0 8320 0 88 84 0 0 4
1133 1124
1133 1199
1370 1199
1370 1178
14 1 95 0 0 8320 0 88 83 0 0 4
1124 1124
1124 1189
1390 1189
1390 1178
1 0 2 0 0 0 0 88 0 0 170 4
1187 1060
1187 1059
1219 1059
1219 1132
9 0 2 0 0 0 0 88 0 0 170 2
1187 1130
1187 1132
10 1 2 0 0 0 0 88 87 0 0 3
1178 1130
1178 1132
1246 1132
2 0 96 0 0 4096 0 88 0 0 172 2
1178 1054
1178 1031
1 3 96 0 0 8320 0 24 88 0 0 4
1694 1033
1694 1031
1169 1031
1169 1054
5 0 41 0 0 0 0 88 0 0 216 3
1151 1060
1151 1036
994 1036
6 0 42 0 0 0 0 88 0 0 215 3
1142 1060
1142 1042
1013 1042
7 0 43 0 0 0 0 88 0 0 214 3
1133 1060
1133 1050
1033 1050
8 0 44 0 0 0 0 88 0 0 213 2
1124 1060
1053 1060
1 10 2 0 0 0 0 89 91 0 0 3
1393 747
1393 745
1363 745
9 0 41 0 0 0 0 90 0 0 216 2
1058 874
994 874
10 0 42 0 0 0 0 90 0 0 215 2
1058 856
1013 856
11 0 43 0 0 0 0 90 0 0 214 2
1058 838
1033 838
12 0 44 0 0 0 0 90 0 0 213 2
1058 820
1053 820
9 1 97 0 0 8320 0 91 29 0 0 4
1354 739
1354 835
1633 835
1633 955
7 1 98 0 0 8320 0 91 28 0 0 4
1336 739
1336 849
1601 849
1601 954
5 1 99 0 0 8320 0 91 27 0 0 4
1318 739
1318 864
1570 864
1570 954
3 1 100 0 0 8320 0 91 26 0 0 4
1300 739
1300 878
1537 878
1537 952
8 1 85 0 0 0 0 91 30 0 0 4
1345 739
1345 918
1386 918
1386 953
6 1 84 0 0 0 0 91 31 0 0 4
1327 739
1327 928
1354 928
1354 952
4 1 83 0 0 4224 0 91 32 0 0 4
1309 739
1309 938
1323 938
1323 952
2 1 82 0 0 8320 0 91 33 0 0 3
1291 739
1290 739
1290 950
1 1 101 0 0 4224 0 34 91 0 0 3
1694 762
1282 762
1282 739
0 7 102 0 0 4096 0 0 92 192 0 3
1129 290
1129 271
1123 271
0 5 102 0 0 0 0 0 92 193 0 3
1129 307
1129 289
1123 289
3 0 102 0 0 0 0 92 0 0 194 3
1123 307
1129 307
1129 325
1 1 102 0 0 4224 0 92 35 0 0 2
1123 325
1686 325
9 0 41 0 0 0 0 92 0 0 216 2
1059 316
994 316
10 0 42 0 0 0 0 92 0 0 215 2
1059 298
1013 298
11 0 43 0 0 0 0 92 0 0 214 2
1059 280
1033 280
12 0 44 0 0 0 0 92 0 0 213 2
1059 262
1053 262
11 2 32 0 0 0 0 94 92 0 0 3
1152 234
1152 316
1123 316
12 4 33 0 0 0 0 94 92 0 0 3
1143 234
1143 298
1123 298
13 6 34 0 0 0 0 94 92 0 0 3
1134 234
1134 280
1123 280
14 8 35 0 0 0 0 94 92 0 0 3
1125 234
1123 234
1123 262
2 0 103 0 0 4096 0 94 0 0 204 2
1179 164
1179 141
1 3 103 0 0 4224 0 36 94 0 0 3
1682 141
1170 141
1170 164
1 0 2 0 0 0 0 94 0 0 207 3
1188 170
1220 170
1220 243
9 0 2 0 0 0 0 94 0 0 207 2
1188 240
1188 243
10 1 2 0 0 0 0 94 93 0 0 3
1179 240
1179 243
1247 243
1 4 3 0 0 4224 0 37 94 0 0 3
112 31
1161 31
1161 170
5 0 41 0 0 0 0 94 0 0 216 3
1152 170
1152 146
994 146
6 0 42 0 0 0 0 94 0 0 215 3
1143 170
1143 152
1013 152
7 0 43 0 0 0 0 94 0 0 214 3
1134 170
1134 160
1033 160
8 0 44 0 0 0 0 94 0 0 213 2
1125 170
1053 170
1 1 44 0 0 4224 0 106 99 0 0 2
1053 112
1053 1225
1 1 43 0 0 4224 0 105 100 0 0 2
1033 112
1033 1225
1 1 42 0 0 4224 0 104 101 0 0 2
1013 112
1013 1225
1 1 41 0 0 4224 0 103 102 0 0 2
994 112
994 1225
1 1 58 0 0 4224 0 107 98 0 0 2
975 112
975 1225
1 1 57 0 0 4224 0 108 97 0 0 2
955 112
955 1225
1 1 56 0 0 4224 0 109 96 0 0 2
935 112
935 1225
1 1 55 0 0 4224 0 110 95 0 0 2
916 112
916 1225
45
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
704 1588 755 1611
717 1598 741 1613
3 HLT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
708 1565 751 1588
721 1575 737 1590
2 JZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1537 757 1560
720 1547 744 1562
3 JMP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1514 757 1537
720 1524 744 1539
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
707 1488 758 1511
720 1498 744 1513
3 MOV
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1460 757 1483
720 1470 744 1485
3 AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
706 1436 757 1459
719 1446 743 1461
3 SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1409 757 1432
720 1419 744 1434
3 ADD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
709 1382 758 1405
721 1392 745 1407
3 LDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 1331 833 1354
803 1341 819 1356
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 1304 829 1327
800 1314 816 1329
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
789 1280 832 1303
802 1290 818 1305
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 1252 833 1275
803 1262 819 1277
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1627 119 1664 143
1638 128 1652 144
2 LA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1653 303 1680 327
1658 307 1674 323
2 EA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1661 739 1694 760
1669 746 1685 761
2 RS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1662 778 1695 799
1670 785 1686 800
2 EB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1653 1027 1690 1051
1663 1035 1679 1051
2 LO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
123 41 160 65
133 49 149 65
2 EP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
121 125 158 149
131 133 147 149
2 LP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
126 338 257 360
135 345 247 361
14 SM  (external)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
119 533 154 555
128 540 144 556
2 CE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
708 78 743 100
717 85 733 101
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
809 364 852 386
818 371 842 387
3 MAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
420 418 527 440
429 425 517 441
11 INPUT & MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
717 667 760 689
726 675 750 691
3 RAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
654 986 689 1008
663 994 679 1010
2 IR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
125 274 162 296
135 281 151 297
2 LM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
130 1058 165 1080
139 1065 155 1081
2 LI
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 1237 168 1259
142 1245 158 1261
2 EI
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
117 7 176 29
126 15 166 31
5 CLOCK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
122 86 157 108
131 93 147 109
2 CP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1647 633 1690 655
1656 640 1680 656
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1758 568 1793 590
1767 575 1783 591
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1791 567 1826 589
1800 575 1816 591
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1822 568 1857 590
1831 575 1847 591
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1725 566 1760 588
1734 574 1750 590
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1645 349 1682 371
1655 356 1671 372
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1275 201 1304 223
1285 208 1293 224
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1373 426 1416 448
1382 434 1406 450
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1409 699 1452 721
1418 706 1442 722
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1163 919 1190 941
1172 926 1180 942
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1504 913 1531 935
1513 920 1521 936
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1229 1051 1304 1073
1238 1058 1294 1074
7 OUT REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1418 1148 1493 1170
1427 1155 1483 1171
7 DISPLAY
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
