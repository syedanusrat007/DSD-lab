CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
80
13 Logic Switch~
5 369 51 0 10 11
0 70 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-7 -20 7 -12
3 V12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
346 0 0
2
42943.7 0
0
13 Logic Switch~
5 337 52 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-7 -20 7 -12
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3169 0 0
2
42943.7 0
0
13 Logic Switch~
5 301 52 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-7 -20 7 -12
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4826 0 0
2
42943.7 0
0
13 Logic Switch~
5 265 51 0 1 11
0 23
0
0 0 21360 782
2 0V
-7 -20 7 -12
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3971 0 0
2
42943.7 0
0
13 Logic Switch~
5 628 53 0 1 11
0 3
0
0 0 21360 782
2 0V
-7 -20 7 -12
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3607 0 0
2
42943.7 0
0
13 Logic Switch~
5 583 51 0 1 11
0 51
0
0 0 21360 782
2 0V
-7 -20 7 -12
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3506 0 0
2
42943.7 0
0
13 Logic Switch~
5 525 53 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-7 -20 7 -12
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7829 0 0
2
42943.7 0
0
13 Logic Switch~
5 481 51 0 1 11
0 26
0
0 0 21360 782
2 0V
-7 -20 7 -12
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3890 0 0
2
42943.7 0
0
13 Logic Switch~
5 170 53 0 1 11
0 67
0
0 0 21360 782
2 0V
-7 -20 7 -12
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3126 0 0
2
42943.7 0
0
13 Logic Switch~
5 117 53 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-7 -20 7 -12
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3935 0 0
2
42943.7 0
0
13 Logic Switch~
5 62 52 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-7 -20 7 -12
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9746 0 0
2
42943.7 0
0
13 Logic Switch~
5 14 55 0 1 11
0 73
0
0 0 21360 782
2 0V
-7 -20 7 -12
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7330 0 0
2
42943.7 0
0
5 4001~
219 982 322 0 3 22
0 3 2 68
0
0 0 624 0
4 4001
-14 -24 14 -16
4 U18D
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 18 0
1 U
3972 0 0
2
42943.8 0
0
5 4001~
219 781 197 0 3 22
0 5 4 72
0
0 0 624 0
4 4001
-14 -24 14 -16
4 U18C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 18 0
1 U
7818 0 0
2
42943.8 0
0
5 4001~
219 705 215 0 3 22
0 6 2 4
0
0 0 624 0
4 4001
-14 -24 14 -16
4 U18B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 18 0
1 U
3818 0 0
2
42943.8 0
0
5 4001~
219 706 182 0 3 22
0 3 7 5
0
0 0 624 0
4 4001
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 18 0
1 U
8835 0 0
2
42943.8 0
0
9 Inverter~
13 76 78 0 2 22
0 7 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U17A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 17 0
1 U
7484 0 0
2
42943.8 0
0
9 2-In AND~
219 1649 312 0 3 22
0 11 10 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
792 0 0
2
42943.7 0
0
9 2-In AND~
219 1658 609 0 3 22
0 13 10 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3826 0 0
2
42943.7 0
0
9 2-In AND~
219 1661 884 0 3 22
0 15 10 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
7958 0 0
2
42943.7 0
0
9 2-In AND~
219 1700 1185 0 3 22
0 16 10 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
6736 0 0
2
42943.7 0
0
9 4-In NOR~
219 2160 112 0 5 22
0 20 19 18 17 21
0
0 0 624 90
4 4002
-14 -24 14 -16
3 U2B
29 -2 50 6
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 2 0
1 U
3755 0 0
2
42943.7 0
0
9 2-In XOR~
219 2048 111 0 3 22
0 8 14 22
0
0 0 624 90
6 74LS86
-21 -24 21 -16
4 U15A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
397 0 0
2
42943.7 0
0
14 Logic Display~
6 2166 62 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5190 0 0
2
42943.7 3
0
14 Logic Display~
6 2110 61 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9188 0 0
2
42943.7 2
0
14 Logic Display~
6 2051 64 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3651 0 0
2
42943.7 1
0
14 Logic Display~
6 2011 64 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3415 0 0
2
42943.7 0
0
14 Logic Display~
6 1689 70 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7597 0 0
2
42943.7 0
0
8 2-In OR~
219 1573 1176 0 3 22
0 29 28 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U13B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
350 0 0
2
42943.7 10
0
9 2-In AND~
219 1490 1167 0 3 22
0 30 14 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
3153 0 0
2
42943.7 9
0
9 2-In AND~
219 1343 1265 0 3 22
0 32 31 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
634 0 0
2
42943.7 8
0
9 2-In XOR~
219 1479 1121 0 3 22
0 30 14 20
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
8956 0 0
2
42943.7 7
0
9 2-In XOR~
219 1383 1112 0 3 22
0 32 31 30
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
3342 0 0
2
42943.7 6
0
8 2-In OR~
219 1157 1162 0 3 22
0 34 33 31
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U13C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
3549 0 0
2
42943.7 5
0
9 2-In AND~
219 1018 1195 0 3 22
0 24 7 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
9177 0 0
2
42943.7 4
0
9 2-In AND~
219 1016 1136 0 3 22
0 26 25 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3387 0 0
2
42943.7 3
0
8 2-In OR~
219 1244 1047 0 3 22
0 35 23 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U13D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
351 0 0
2
42943.7 2
0
9 2-In AND~
219 1121 1038 0 3 22
0 27 36 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
3127 0 0
2
42943.7 1
0
9 2-In XOR~
219 1006 1079 0 3 22
0 26 7 36
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
559 0 0
2
42943.7 0
0
14 Logic Display~
6 1729 70 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8488 0 0
2
42943.7 0
0
8 2-In OR~
219 1565 875 0 3 22
0 41 40 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
3392 0 0
2
42943.7 10
0
9 2-In AND~
219 1482 866 0 3 22
0 42 12 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3952 0 0
2
42943.7 9
0
9 2-In AND~
219 1335 964 0 3 22
0 44 43 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
8186 0 0
2
42943.7 8
0
9 2-In XOR~
219 1471 820 0 3 22
0 42 12 19
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
6571 0 0
2
42943.7 7
0
9 2-In XOR~
219 1375 811 0 3 22
0 44 43 42
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
6167 0 0
2
42943.7 6
0
8 2-In OR~
219 1149 861 0 3 22
0 46 45 43
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3566 0 0
2
42943.7 5
0
9 2-In AND~
219 1010 894 0 3 22
0 38 7 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3371 0 0
2
42943.7 4
0
9 2-In AND~
219 1008 835 0 3 22
0 39 25 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
4395 0 0
2
42943.7 3
0
8 2-In OR~
219 1236 746 0 3 22
0 47 37 44
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
6822 0 0
2
42943.7 2
0
9 2-In AND~
219 1113 737 0 3 22
0 27 48 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
8953 0 0
2
42943.7 1
0
9 2-In XOR~
219 998 778 0 3 22
0 39 7 48
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
4635 0 0
2
42943.7 0
0
14 Logic Display~
6 1788 67 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6596 0 0
2
42943.7 0
0
9 2-In XOR~
219 998 503 0 3 22
0 51 7 60
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3813 0 0
2
42943.7 11
0
9 2-In AND~
219 1113 462 0 3 22
0 27 60 59
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
5639 0 0
2
42943.7 10
0
8 2-In OR~
219 1236 471 0 3 22
0 59 49 56
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
429 0 0
2
42943.7 9
0
9 2-In AND~
219 1008 560 0 3 22
0 51 25 58
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
5832 0 0
2
42943.7 8
0
9 2-In AND~
219 1010 619 0 3 22
0 50 7 57
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
8856 0 0
2
42943.7 7
0
8 2-In OR~
219 1149 586 0 3 22
0 58 57 55
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
469 0 0
2
42943.7 6
0
9 2-In XOR~
219 1375 536 0 3 22
0 56 55 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
4529 0 0
2
42943.7 4
0
9 2-In XOR~
219 1471 545 0 3 22
0 54 9 18
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
88 0 0
2
42943.7 3
0
9 2-In AND~
219 1335 689 0 3 22
0 56 55 52
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3894 0 0
2
42943.7 2
0
9 2-In AND~
219 1482 591 0 3 22
0 54 9 53
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
6890 0 0
2
42943.7 1
0
8 2-In OR~
219 1565 600 0 3 22
0 53 52 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3257 0 0
2
42943.7 0
0
14 Logic Display~
6 1844 68 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6612 0 0
2
42943.7 0
0
8 2-In OR~
219 1554 303 0 3 22
0 62 61 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3556 0 0
2
42943.7 0
0
9 2-In AND~
219 1471 294 0 3 22
0 64 63 62
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9143 0 0
2
42943.7 0
0
9 2-In AND~
219 1324 392 0 3 22
0 66 65 61
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8186 0 0
2
42943.7 0
0
9 2-In XOR~
219 1460 248 0 3 22
0 64 63 17
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3754 0 0
2
42943.7 0
0
9 2-In XOR~
219 1364 239 0 3 22
0 66 65 64
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8708 0 0
2
42943.7 0
0
9 2-In AND~
219 1145 364 0 3 22
0 10 67 63
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3338 0 0
2
42943.7 0
0
8 2-In OR~
219 1138 289 0 3 22
0 69 68 65
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5546 0 0
2
42943.7 0
0
9 2-In AND~
219 997 263 0 3 22
0 3 25 69
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3295 0 0
2
42943.7 0
0
8 2-In OR~
219 1225 174 0 3 22
0 71 70 66
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4923 0 0
2
42943.7 0
0
9 2-In AND~
219 1102 165 0 3 22
0 27 72 71
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3248 0 0
2
42943.7 0
0
9 4-In NOR~
219 816 156 0 5 22
0 10 25 74 75 27
0
0 0 624 0
4 4002
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 1 2 0
1 U
3139 0 0
2
42943.7 0
0
9 Inverter~
13 644 74 0 2 22
0 3 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3285 0 0
2
42943.7 0
0
9 Inverter~
13 597 74 0 2 22
0 51 50
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
336 0 0
2
42943.7 0
0
9 Inverter~
13 539 74 0 2 22
0 39 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6582 0 0
2
42943.7 0
0
9 Inverter~
13 496 73 0 2 22
0 26 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3546 0 0
2
42943.7 0
0
9 Inverter~
13 30 78 0 2 22
0 73 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
893 0 0
2
42943.7 0
0
142
2 0 2 0 0 4096 0 13 0 0 9 2
969 331
97 331
1 0 3 0 0 4096 0 13 0 0 135 2
969 313
628 313
3 2 4 0 0 4224 0 15 14 0 0 4
744 215
759 215
759 206
768 206
3 1 5 0 0 4224 0 16 14 0 0 4
745 182
760 182
760 188
768 188
2 0 2 0 0 0 0 15 0 0 9 2
692 224
97 224
1 0 6 0 0 4096 0 15 0 0 121 2
692 206
665 206
2 0 7 0 0 4096 0 16 0 0 141 2
693 191
62 191
1 0 3 0 0 0 0 16 0 0 135 2
693 173
628 173
2 0 2 0 0 4224 0 17 0 0 0 2
97 78
97 1361
1 0 7 0 0 0 0 17 0 0 141 2
61 78
62 78
1 0 8 0 0 8192 0 23 0 0 25 3
2042 130
2042 138
2011 138
2 0 9 0 0 4096 0 60 0 0 13 2
1455 554
1427 554
3 2 9 0 0 12416 0 18 62 0 0 6
1670 312
1682 312
1682 484
1427 484
1427 600
1458 600
2 0 10 0 0 12288 0 18 0 0 110 5
1625 321
1595 321
1595 410
739 410
739 355
3 1 11 0 0 4224 0 65 18 0 0 2
1587 303
1625 303
2 0 10 0 0 12288 0 19 0 0 125 4
1634 618
1599 618
1599 645
51 645
2 0 10 0 0 12288 0 20 0 0 125 4
1637 893
1601 893
1601 929
51 929
2 0 10 0 0 12416 0 21 0 0 125 4
1676 1194
1624 1194
1624 1224
51 1224
2 0 12 0 0 4096 0 44 0 0 20 2
1455 829
1426 829
3 2 12 0 0 8320 0 19 42 0 0 5
1679 609
1679 747
1426 747
1426 875
1458 875
3 1 13 0 0 4224 0 63 19 0 0 2
1598 600
1634 600
2 0 14 0 0 4096 0 32 0 0 23 2
1463 1130
1437 1130
2 0 14 0 0 12288 0 30 0 0 33 5
1466 1176
1437 1176
1437 991
1767 991
1767 898
3 1 15 0 0 4224 0 41 20 0 0 2
1598 875
1637 875
1 3 8 0 0 4224 0 27 21 0 0 3
2011 82
2011 1185
1721 1185
3 1 16 0 0 4224 0 29 21 0 0 2
1606 1176
1676 1176
4 0 17 0 0 8192 0 22 0 0 104 3
2180 135
2180 172
1844 172
3 0 18 0 0 8192 0 22 0 0 78 3
2171 135
2171 163
1788 163
2 0 19 0 0 8192 0 22 0 0 64 3
2162 135
2162 147
1729 147
1 0 20 0 0 4096 0 22 0 0 32 2
2153 135
2110 135
5 1 21 0 0 4224 0 22 24 0 0 2
2166 79
2166 80
1 0 20 0 0 8192 0 25 0 0 43 3
2110 79
2110 178
1689 178
2 3 14 0 0 4224 0 23 20 0 0 5
2060 130
2060 898
1714 898
1714 884
1682 884
3 1 22 0 0 4224 0 23 26 0 0 2
2051 81
2051 82
2 0 23 0 0 12288 0 37 0 0 134 4
1231 1056
1154 1056
1154 1106
265 1106
2 0 7 0 0 4096 0 35 0 0 141 2
994 1204
62 1204
1 0 24 0 0 4096 0 35 0 0 124 2
994 1186
517 1186
2 0 25 0 0 4096 0 36 0 0 140 2
992 1145
117 1145
1 0 26 0 0 4096 0 36 0 0 138 2
992 1127
481 1127
2 0 7 0 0 0 0 39 0 0 141 2
990 1088
62 1088
1 0 26 0 0 0 0 39 0 0 138 2
990 1070
481 1070
0 1 27 0 0 4224 0 0 38 118 0 3
933 156
933 1029
1097 1029
3 1 20 0 0 8320 0 32 28 0 0 3
1512 1121
1689 1121
1689 88
3 2 28 0 0 4224 0 31 29 0 0 4
1364 1265
1537 1265
1537 1185
1560 1185
3 1 29 0 0 4224 0 30 29 0 0 2
1511 1167
1560 1167
1 0 30 0 0 8192 0 30 0 0 49 3
1466 1158
1452 1158
1452 1112
2 0 31 0 0 8192 0 31 0 0 50 3
1319 1274
1264 1274
1264 1162
1 0 32 0 0 8320 0 31 0 0 51 3
1319 1256
1304 1256
1304 1047
3 1 30 0 0 4224 0 33 32 0 0 2
1416 1112
1463 1112
3 2 31 0 0 4224 0 34 33 0 0 4
1190 1162
1356 1162
1356 1121
1367 1121
3 1 32 0 0 0 0 37 33 0 0 4
1277 1047
1355 1047
1355 1103
1367 1103
3 2 33 0 0 4224 0 35 34 0 0 4
1039 1195
1126 1195
1126 1171
1144 1171
3 1 34 0 0 4224 0 36 34 0 0 4
1037 1136
1126 1136
1126 1153
1144 1153
3 1 35 0 0 4224 0 38 37 0 0 2
1142 1038
1231 1038
3 2 36 0 0 4224 0 39 38 0 0 4
1039 1079
1078 1079
1078 1047
1097 1047
2 0 37 0 0 12288 0 49 0 0 133 4
1223 755
1153 755
1153 807
301 807
2 0 7 0 0 0 0 47 0 0 141 2
986 903
62 903
1 0 38 0 0 4096 0 47 0 0 123 2
986 885
560 885
2 0 25 0 0 0 0 48 0 0 140 2
984 844
117 844
1 0 39 0 0 4096 0 48 0 0 137 2
984 826
525 826
2 0 7 0 0 0 0 51 0 0 141 2
982 787
62 787
1 0 39 0 0 0 0 51 0 0 137 2
982 769
525 769
0 1 27 0 0 0 0 0 50 118 0 3
957 156
957 728
1089 728
3 1 19 0 0 8320 0 44 40 0 0 3
1504 820
1729 820
1729 88
3 2 40 0 0 4224 0 43 41 0 0 4
1356 964
1529 964
1529 884
1552 884
3 1 41 0 0 4224 0 42 41 0 0 2
1503 866
1552 866
1 0 42 0 0 8192 0 42 0 0 70 3
1458 857
1444 857
1444 811
2 0 43 0 0 8192 0 43 0 0 71 3
1311 973
1256 973
1256 861
1 0 44 0 0 8320 0 43 0 0 72 3
1311 955
1296 955
1296 746
3 1 42 0 0 4224 0 45 44 0 0 2
1408 811
1455 811
3 2 43 0 0 4224 0 46 45 0 0 4
1182 861
1348 861
1348 820
1359 820
3 1 44 0 0 0 0 49 45 0 0 4
1269 746
1347 746
1347 802
1359 802
3 2 45 0 0 4224 0 47 46 0 0 4
1031 894
1118 894
1118 870
1136 870
3 1 46 0 0 4224 0 48 46 0 0 4
1029 835
1118 835
1118 852
1136 852
3 1 47 0 0 4224 0 50 49 0 0 2
1134 737
1223 737
3 2 48 0 0 4224 0 51 50 0 0 4
1031 778
1070 778
1070 746
1089 746
2 0 49 0 0 12288 0 55 0 0 132 4
1223 480
1140 480
1140 528
337 528
3 1 18 0 0 8320 0 60 52 0 0 3
1504 545
1788 545
1788 85
2 0 7 0 0 0 0 57 0 0 141 2
986 628
62 628
1 0 50 0 0 4096 0 57 0 0 122 2
986 610
618 610
2 0 25 0 0 0 0 56 0 0 140 2
984 569
117 569
1 0 51 0 0 4096 0 56 0 0 136 2
984 551
583 551
2 0 7 0 0 0 0 53 0 0 141 2
982 512
62 512
1 0 51 0 0 0 0 53 0 0 136 2
982 494
583 494
0 1 27 0 0 0 0 0 54 118 0 3
1046 156
1046 453
1089 453
3 2 52 0 0 4224 0 61 63 0 0 4
1356 689
1529 689
1529 609
1552 609
3 1 53 0 0 4224 0 62 63 0 0 2
1503 591
1552 591
1 0 54 0 0 8192 0 62 0 0 91 3
1458 582
1444 582
1444 536
2 0 55 0 0 8192 0 61 0 0 92 3
1311 698
1256 698
1256 586
1 0 56 0 0 8320 0 61 0 0 93 3
1311 680
1296 680
1296 471
3 1 54 0 0 4224 0 59 60 0 0 2
1408 536
1455 536
3 2 55 0 0 4224 0 58 59 0 0 4
1182 586
1348 586
1348 545
1359 545
3 1 56 0 0 0 0 55 59 0 0 4
1269 471
1347 471
1347 527
1359 527
3 2 57 0 0 4224 0 57 58 0 0 4
1031 619
1118 619
1118 595
1136 595
3 1 58 0 0 4224 0 56 58 0 0 4
1029 560
1118 560
1118 577
1136 577
3 1 59 0 0 4224 0 54 55 0 0 2
1134 462
1223 462
3 2 60 0 0 4224 0 53 54 0 0 4
1031 503
1070 503
1070 471
1089 471
3 2 61 0 0 4224 0 67 65 0 0 4
1345 392
1518 392
1518 312
1541 312
3 1 62 0 0 4224 0 66 65 0 0 2
1492 294
1541 294
2 0 63 0 0 4096 0 66 0 0 105 2
1447 303
1412 303
1 0 64 0 0 8192 0 66 0 0 106 3
1447 285
1433 285
1433 239
2 0 65 0 0 8192 0 67 0 0 107 3
1300 401
1245 401
1245 289
1 0 66 0 0 8320 0 67 0 0 108 3
1300 383
1285 383
1285 174
3 1 17 0 0 4224 0 68 64 0 0 3
1493 248
1844 248
1844 86
3 2 63 0 0 4224 0 70 68 0 0 4
1166 364
1412 364
1412 257
1444 257
3 1 64 0 0 4224 0 69 68 0 0 2
1397 239
1444 239
3 2 65 0 0 4224 0 71 69 0 0 4
1171 289
1337 289
1337 248
1348 248
3 1 66 0 0 0 0 73 69 0 0 4
1258 174
1336 174
1336 230
1348 230
2 0 67 0 0 4096 0 70 0 0 139 2
1121 373
170 373
1 0 10 0 0 0 0 70 0 0 125 2
1121 355
51 355
3 2 68 0 0 4224 0 13 71 0 0 4
1021 322
1107 322
1107 298
1125 298
3 1 69 0 0 4224 0 72 71 0 0 4
1018 263
1107 263
1107 280
1125 280
2 0 25 0 0 0 0 72 0 0 140 2
973 272
117 272
1 0 3 0 0 4096 0 72 0 0 135 2
973 254
628 254
2 0 70 0 0 12288 0 73 0 0 131 4
1212 183
1124 183
1124 234
369 234
3 1 71 0 0 4224 0 74 73 0 0 2
1123 165
1212 165
3 2 72 0 0 4224 0 14 74 0 0 6
820 197
1010 197
1010 206
1059 206
1059 174
1078 174
5 1 27 0 0 0 0 75 74 0 0 2
855 156
1078 156
2 0 25 0 0 0 0 75 0 0 140 2
799 152
117 152
1 0 10 0 0 0 0 75 0 0 125 2
799 143
51 143
2 0 6 0 0 4224 0 76 0 0 0 2
665 74
665 1359
2 0 50 0 0 4224 0 77 0 0 0 2
618 74
618 1357
2 0 38 0 0 4224 0 78 0 0 0 2
560 74
560 1361
2 0 24 0 0 4224 0 79 0 0 0 2
517 73
517 1359
2 0 10 0 0 128 0 80 0 0 0 2
51 78
51 1354
1 0 3 0 0 0 0 76 0 0 135 2
629 74
628 74
1 0 51 0 0 0 0 77 0 0 136 2
582 74
583 74
1 0 39 0 0 0 0 78 0 0 137 2
524 74
525 74
1 0 26 0 0 0 0 79 0 0 138 2
481 73
481 73
1 0 73 0 0 4096 0 80 0 0 142 2
15 78
14 78
1 0 70 0 0 4224 0 1 0 0 0 2
369 63
369 1354
1 0 49 0 0 4224 0 2 0 0 0 2
337 64
337 1353
1 0 37 0 0 4224 0 3 0 0 0 2
301 64
301 1347
1 0 23 0 0 4224 0 4 0 0 0 2
265 63
265 1349
1 0 3 0 0 4224 0 5 0 0 0 2
628 65
628 1358
1 0 51 0 0 4224 0 6 0 0 0 2
583 63
583 1355
1 0 39 0 0 4224 0 7 0 0 0 2
525 65
525 1358
1 0 26 0 0 4224 0 8 0 0 0 2
481 63
481 1355
1 0 67 0 0 4224 0 9 0 0 0 2
170 65
170 1352
1 0 25 0 0 4224 0 10 0 0 0 2
117 65
117 1352
1 0 7 0 0 4224 0 11 0 0 0 2
62 64
62 1349
1 0 73 0 0 4224 0 12 0 0 0 2
14 67
14 1350
47
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 33
345 190 664 221
352 194 656 215
33 (B1+S1)' nor (B1'+S1')'=B1 xor S1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 15
711 285 872 316
718 289 864 310
15 (B1+S1')'=B1'S1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 50
877 8 966 143
884 12 958 117
50 and ic-6
or ic -3
xor ic-3
not ic -1
nor ic -2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1079 149 1119 180
1086 153 1111 174
2 24
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1544 290 1581 321
1551 294 1573 315
2 12
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
2034 91 2071 122
2041 95 2063 116
2 12
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
2154 95 2182 126
2161 99 2174 120
1 2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
977 308 1004 339
984 312 996 333
1 4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
637 80 664 111
644 84 656 105
1 6
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 15
696 101 867 132
703 105 859 126
15 (S2'+S0)'=S2S0'
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
2152 12 2181 43
2159 16 2173 37
1 Z
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
2096 11 2123 42
2103 15 2115 36
1 S
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
2038 14 2066 45
2045 18 2058 39
1 V
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1992 14 2021 45
1999 18 2013 39
1 C
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1668 15 1709 46
1675 19 1701 40
2 F4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1563 1124 1604 1155
1570 1128 1596 1149
2 C5
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1459 1056 1500 1087
1466 1060 1492 1081
2 F4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1152 1112 1186 1143
1156 1116 1181 1137
2 Y4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1229 988 1263 1019
1233 992 1258 1013
2 X4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1555 823 1596 854
1562 827 1588 848
2 C4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1555 548 1596 579
1562 552 1588 573
2 C3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1544 251 1586 282
1551 255 1578 276
2 C2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1708 13 1749 44
1715 17 1741 38
2 F3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1144 811 1178 842
1148 815 1173 836
2 Y3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1204 693 1238 724
1208 697 1233 718
2 X3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1451 755 1492 786
1458 759 1484 780
2 F3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1769 13 1811 44
1776 17 1803 38
2 F2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1451 480 1493 511
1458 484 1485 505
2 F2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1144 536 1179 567
1148 540 1174 561
2 Y2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1204 418 1239 449
1208 422 1234 443
2 X2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1826 12 1864 43
1833 16 1856 37
2 F1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1440 183 1478 214
1447 187 1470 208
2 F1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1122 317 1160 348
1129 321 1152 342
2 Z1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1133 239 1170 270
1140 243 1162 264
2 Y1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1193 121 1230 152
1200 125 1222 146
2 X1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
613 -4 646 27
617 0 641 21
2 B1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
562 -4 599 27
566 0 594 21
2 B2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
508 -4 544 27
512 0 539 21
2 B3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
461 -4 497 27
465 0 492 21
2 B4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
356 -4 387 27
360 0 382 21
2 A1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
323 -4 358 27
327 0 353 21
2 A2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
288 -4 322 27
292 0 317 21
2 A3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
250 -4 284 27
254 0 279 21
2 A4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
152 -4 192 27
156 0 187 21
3 Cin
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
103 -4 137 27
107 0 132 21
2 S0
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
48 -4 78 27
52 0 73 21
2 S1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
-2 -3 32 28
2 1 27 22
2 S2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
