CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
280 1940 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
30 C:\Program Files (x86)\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
137
13 Logic Switch~
5 322 1720 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 180
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89815e-315 0
0
13 Logic Switch~
5 1542 1101 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89815e-315 0
0
13 Logic Switch~
5 1509 1101 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89815e-315 5.26354e-315
0
13 Logic Switch~
5 1472 1101 0 1 11
0 41
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89815e-315 5.30499e-315
0
13 Logic Switch~
5 1437 1099 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89815e-315 5.32571e-315
0
13 Logic Switch~
5 1216 1098 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89815e-315 5.34643e-315
0
13 Logic Switch~
5 1176 1096 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89815e-315 5.3568e-315
0
13 Logic Switch~
5 1138 1096 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.89815e-315 5.36716e-315
0
13 Logic Switch~
5 1101 1095 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.89815e-315 5.37752e-315
0
13 Logic Switch~
5 264 766 0 10 11
0 78 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.89815e-315 5.38788e-315
0
13 Logic Switch~
5 233 745 0 10 11
0 79 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-1 -15 13 -7
2 V7
2 -26 16 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.89815e-315 5.39306e-315
0
13 Logic Switch~
5 201 724 0 1 11
0 80
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.89815e-315 5.39824e-315
0
13 Logic Switch~
5 188 688 0 1 11
0 77
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
5.89815e-315 5.40342e-315
0
13 Logic Switch~
5 201 600 0 10 11
0 81 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.89815e-315 5.4086e-315
0
14 Logic Display~
6 1529 2532 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L61
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
42987.8 0
0
14 Logic Display~
6 1423 2537 0 1 2
10 4
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L60
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
42987.8 0
0
5 4071~
219 1443 2285 0 3 22
0 3 4 5
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U6B
32 -7 53 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
5616 0 0
2
42987.8 0
0
14 Logic Display~
6 382 1628 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L59
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89815e-315 0
0
7 Pulser~
4 337 1654 0 10 12
0 111 112 7 113 0 0 5 5 6
7
0
0 0 4656 0
0
3 V17
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
317 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1342 498 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L58
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89815e-315 5.41896e-315
0
14 Logic Display~
6 1310 498 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L57
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.89815e-315 5.42414e-315
0
14 Logic Display~
6 1277 500 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L56
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89815e-315 5.42933e-315
0
14 Logic Display~
6 1246 502 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L55
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89815e-315 5.43192e-315
0
14 Logic Display~
6 1529 412 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L54
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89815e-315 5.43451e-315
0
14 Logic Display~
6 1484 1374 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L53
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89815e-315 5.4371e-315
0
14 Logic Display~
6 1461 1378 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L52
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89815e-315 5.43969e-315
0
14 Logic Display~
6 1431 1379 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L51
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89815e-315 5.44228e-315
0
14 Logic Display~
6 1403 1378 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L50
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89815e-315 5.44487e-315
0
7 Ground~
168 1329 1426 0 1 3
0 2
0
0 0 53360 512
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
961 0 0
2
5.89815e-315 5.44746e-315
0
7 74LS173
129 1236 1366 0 14 29
0 24 25 25 8 30 31 32 33 24
24 26 27 28 29
0
0 0 4848 270
7 74LS173
-24 -51 25 -43
3 U32
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3178 0 0
2
5.89815e-315 5.45005e-315
0
7 Ground~
168 1450 876 0 1 3
0 2
0
0 0 53360 782
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
5.89815e-315 5.45264e-315
0
9 Inverter~
13 1375 2275 0 2 22
0 3 43
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U12F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
3951 0 0
2
5.89815e-315 5.45523e-315
0
7 74LS126
116 1060 928 0 12 25
0 34 35 34 36 34 37 34 38 30
31 32 33
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
3 U31
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
8885 0 0
2
5.89815e-315 5.45782e-315
0
7 74LS257
147 1321 840 0 14 29
0 43 35 42 36 41 37 40 38 39
2 44 45 46 47
0
0 0 4848 90
7 74LS257
-24 -60 25 -52
3 U30
53 -6 74 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3780 0 0
2
5.89815e-315 5.46041e-315
0
7 74LS181
132 1232 651 0 22 45
0 48 4 5 6 49 50 51 52 44
45 46 47 6 3 114 115 116 117 22
21 20 19
0
0 0 4848 180
7 74LS181
-24 -69 25 -61
3 U29
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
9265 0 0
2
5.89815e-315 5.463e-315
0
7 74LS126
116 1091 630 0 12 25
0 53 22 53 21 53 20 53 19 30
31 32 33
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
3 U28
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
9442 0 0
2
5.89815e-315 5.46559e-315
0
14 Logic Display~
6 1321 194 0 1 2
10 52
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L49
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89815e-315 5.46818e-315
0
14 Logic Display~
6 1371 200 0 1 2
10 51
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L48
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89815e-315 5.47077e-315
0
14 Logic Display~
6 1416 203 0 1 2
10 50
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L47
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89815e-315 5.47207e-315
0
14 Logic Display~
6 1438 202 0 1 2
10 49
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L46
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89815e-315 5.47336e-315
0
9 4-In NOR~
219 1461 430 0 5 22
0 52 51 50 49 23
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U27A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 15 0
1 U
7168 0 0
2
5.89815e-315 5.47466e-315
0
7 Ground~
168 1282 301 0 1 3
0 2
0
0 0 53360 782
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
5.89815e-315 5.47595e-315
0
7 74LS126
116 1079 418 0 12 25
0 54 49 54 50 54 51 54 52 30
31 32 33
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
3 U26
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
4139 0 0
2
5.89815e-315 5.47725e-315
0
7 74LS173
129 1164 298 0 14 29
0 2 55 55 8 30 31 32 33 2
2 49 50 51 52
0
0 0 4848 270
7 74LS173
-24 -51 25 -43
3 U25
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6435 0 0
2
5.89815e-315 5.47854e-315
0
14 Logic Display~
6 1004 1671 0 1 2
10 33
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L45
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.89815e-315 5.47984e-315
0
14 Logic Display~
6 961 1668 0 1 2
10 32
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L44
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
5.89815e-315 5.48113e-315
0
14 Logic Display~
6 922 1665 0 1 2
10 31
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L43
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.89815e-315 5.48243e-315
0
14 Logic Display~
6 886 1663 0 1 2
10 30
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L42
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.89815e-315 5.48372e-315
0
14 Logic Display~
6 846 1664 0 1 2
10 67
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L41
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.89815e-315 5.48502e-315
0
14 Logic Display~
6 807 1663 0 1 2
10 68
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.89815e-315 5.48631e-315
0
14 Logic Display~
6 769 1662 0 1 2
10 69
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L39
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.89815e-315 5.48761e-315
0
14 Logic Display~
6 737 1670 0 1 2
10 70
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L38
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.89815e-315 5.4889e-315
0
7 Ground~
168 457 1666 0 1 3
0 2
0
0 0 53360 512
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6118 0 0
2
5.89815e-315 5.4902e-315
0
9 2-In XOR~
219 463 1642 0 3 22
0 2 60 61
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U24A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
34 0 0
2
5.89815e-315 5.49149e-315
0
7 Ground~
168 663 1348 0 1 3
0 2
0
0 0 53360 512
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
5.89815e-315 5.49279e-315
0
7 74LS126
116 662 1449 0 12 25
0 62 66 62 65 62 64 62 63 33
32 31 30
0
0 0 4848 0
7 74LS126
-24 -51 25 -43
3 U23
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
319 0 0
2
5.89815e-315 5.49408e-315
0
7 74LS173
129 544 1292 0 14 29
0 2 71 71 8 33 32 31 30 2
2 66 65 64 63
0
0 0 4848 270
7 74LS173
-24 -51 25 -43
3 U22
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3976 0 0
2
5.89815e-315 5.49538e-315
0
7 74LS173
129 337 1292 0 14 29
0 61 71 71 8 67 68 69 118 2
2 59 58 57 56
0
0 0 4848 270
7 74LS173
-24 -51 25 -43
3 U21
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
7634 0 0
2
5.89815e-315 5.49667e-315
0
7 Ground~
168 365 952 0 1 3
0 2
0
0 0 53360 602
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
523 0 0
2
5.89815e-315 5.49797e-315
0
6 PROM32
80 602 953 0 14 29
0 72 2 73 74 75 76 70 69 68
67 30 31 32 33
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U20
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
6748 0 0
2
5.89815e-315 5.49926e-315
0
BKGACAAAAAAAAAAAAAAAAFAAAAAAAAAFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 Ground~
168 371 735 0 1 3
0 2
0
0 0 53360 602
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6901 0 0
2
5.89815e-315 5.50056e-315
0
7 Ground~
168 692 586 0 1 3
0 2
0
0 0 53360 782
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
842 0 0
2
5.89815e-315 5.50185e-315
0
7 74LS257
147 457 797 0 14 29
0 81 82 78 83 79 84 80 85 77
2 76 75 74 73
0
0 0 4848 270
7 74LS257
-24 -60 25 -52
3 U19
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3277 0 0
2
5.89815e-315 5.50315e-315
0
7 74LS173
129 571 597 0 14 29
0 2 86 86 8 33 32 31 30 2
2 82 83 84 85
0
0 0 4848 270
7 74LS173
-24 -51 25 -43
3 U18
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4212 0 0
2
5.89815e-315 5.50444e-315
0
7 Ground~
168 339 172 0 1 3
0 2
0
0 0 53360 692
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4720 0 0
2
5.89815e-315 5.50574e-315
0
2 +V
167 364 169 0 1 3
0 89
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5551 0 0
2
5.89815e-315 5.50703e-315
0
7 74LS154
95 242 1904 0 22 45
0 2 2 56 57 58 59 119 120 121
122 123 124 10 11 12 13 14 15 16
17 18 125
0
0 0 4848 270
7 74LS154
-24 -87 25 -79
3 U15
81 -2 102 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
6986 0 0
2
5.89815e-315 5.50833e-315
0
7 74LS164
127 412 1860 0 12 25
0 105 105 8 106 126 127 128 129 93
9 88 60
0
0 0 4848 0
7 74LS164
-24 -51 25 -43
3 U14
-10 -52 11 -44
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
8745 0 0
2
5.89815e-315 5.50963e-315
0
2 +V
167 348 1883 0 1 3
0 106
0
0 0 54256 90
3 10V
-1 -13 20 -5
2 V1
1 -21 15 -13
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9592 0 0
2
5.89815e-315 5.51092e-315
0
9 3-In NOR~
219 317 1825 0 4 22
0 60 88 9 105
0
0 0 624 0
6 74LS27
-21 -24 21 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 13 0
1 U
8748 0 0
2
5.89815e-315 5.51222e-315
0
7 Ground~
168 287 1867 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
5.89815e-315 5.51286e-315
0
9 Inverter~
13 347 1974 0 2 22
0 18 100
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
631 0 0
2
5.89815e-315 5.51351e-315
0
9 Inverter~
13 347 2010 0 2 22
0 17 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
9466 0 0
2
5.89815e-315 5.51416e-315
0
9 Inverter~
13 347 2048 0 2 22
0 16 3
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
3266 0 0
2
5.89815e-315 5.51481e-315
0
9 Inverter~
13 345 2078 0 2 22
0 15 4
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
7693 0 0
2
5.89815e-315 5.51545e-315
0
9 Inverter~
13 343 2108 0 2 22
0 14 94
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
3723 0 0
2
5.89815e-315 5.5161e-315
0
9 Inverter~
13 343 2136 0 2 22
0 13 96
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
3440 0 0
2
5.89815e-315 5.51675e-315
0
9 Inverter~
13 343 2158 0 2 22
0 12 101
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
6263 0 0
2
5.89815e-315 5.5174e-315
0
9 Inverter~
13 341 2189 0 2 22
0 11 103
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
4900 0 0
2
5.89815e-315 5.51804e-315
0
9 Inverter~
13 342 2214 0 2 22
0 10 104
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
8783 0 0
2
5.89815e-315 5.51869e-315
0
14 Logic Display~
6 387 2479 0 1 2
10 60
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
5.89815e-315 5.51934e-315
0
14 Logic Display~
6 428 2494 0 1 2
10 88
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3215 0 0
2
5.89815e-315 5.51999e-315
0
9 2-In AND~
219 513 2249 0 3 22
0 23 103 102
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U9D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
7903 0 0
2
5.89815e-315 5.52063e-315
0
8 2-In OR~
219 497 2306 0 3 22
0 101 102 90
0
0 0 624 782
5 74F32
-18 -24 17 -16
3 U3B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7121 0 0
2
5.89815e-315 5.52128e-315
0
5 4011~
219 492 2399 0 3 22
0 90 9 87
0
0 0 624 270
4 4011
-7 -24 21 -16
4 U11B
16 -7 44 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 11 0
1 U
4484 0 0
2
5.89815e-315 5.52193e-315
0
14 Logic Display~
6 493 2472 0 1 2
10 87
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.89815e-315 5.52258e-315
0
9 2-In AND~
219 638 2250 0 3 22
0 100 9 91
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U9C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
7804 0 0
2
5.89815e-315 5.52322e-315
0
9 2-In AND~
219 732 2254 0 3 22
0 100 93 97
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U9B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
5523 0 0
2
5.89815e-315 5.52387e-315
0
5 4001~
219 715 2318 0 3 22
0 97 88 72
0
0 0 624 270
4 4001
-14 -24 14 -16
3 U8B
31 -10 52 -2
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 8 0
1 U
3330 0 0
2
5.89815e-315 5.52452e-315
0
14 Logic Display~
6 627 2488 0 1 2
10 86
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
5.89815e-315 5.52517e-315
0
14 Logic Display~
6 721 2481 0 1 2
10 72
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
5.89815e-315 5.52581e-315
0
9 Inverter~
13 784 2372 0 2 22
0 130 71
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U4B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 2 4 0
1 U
3685 0 0
2
5.89815e-315 5.52646e-315
0
14 Logic Display~
6 786 2481 0 1 2
10 71
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
5.89815e-315 5.52711e-315
0
5 4011~
219 817 2302 0 3 22
0 100 9 62
0
0 0 624 270
4 4011
-7 -24 21 -16
4 U11A
16 -7 44 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 11 0
1 U
6343 0 0
2
5.89815e-315 5.52776e-315
0
14 Logic Display~
6 836 2484 0 1 2
10 62
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
5.89815e-315 5.52841e-315
0
8 4-In OR~
219 905 2254 0 5 22
0 6 3 4 94 99
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U10A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
9156 0 0
2
5.89815e-315 5.52905e-315
0
9 2-In AND~
219 901 2318 0 3 22
0 99 9 98
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U9A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5776 0 0
2
5.89815e-315 5.5297e-315
0
5 4001~
219 890 2384 0 3 22
0 98 97 55
0
0 0 624 270
4 4001
-14 -24 14 -16
3 U8A
31 -10 52 -2
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 8 0
1 U
7207 0 0
2
5.89815e-315 5.53035e-315
0
14 Logic Display~
6 895 2489 0 1 2
10 55
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
5.89815e-315 5.531e-315
0
9 2-In AND~
219 982 2260 0 3 22
0 96 9 54
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U5D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3760 0 0
2
5.89815e-315 5.53164e-315
0
14 Logic Display~
6 980 2481 0 1 2
10 54
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
5.89815e-315 5.53229e-315
0
8 3-In OR~
219 1052 2258 0 4 22
0 6 3 4 95
0
0 0 624 270
4 4075
-14 -24 14 -16
3 U7A
32 -7 53 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
9767 0 0
2
5.89815e-315 5.53294e-315
0
9 2-In AND~
219 1049 2330 0 3 22
0 95 9 53
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U5C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7978 0 0
2
5.89815e-315 5.53359e-315
0
14 Logic Display~
6 1047 2491 0 1 2
10 53
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L10
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3142 0 0
2
5.89815e-315 5.53423e-315
0
14 Logic Display~
6 1150 2481 0 1 2
10 3
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L11
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
5.89815e-315 5.53553e-315
0
5 4071~
219 1194 2260 0 3 22
0 6 3 48
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U6A
32 -7 53 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
659 0 0
2
5.89815e-315 5.53618e-315
0
14 Logic Display~
6 1209 2497 0 1 2
10 48
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L12
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
5.89815e-315 5.53682e-315
0
9 2-In AND~
219 1331 2272 0 3 22
0 94 9 34
0
0 0 624 270
5 74F08
-18 -24 17 -16
3 U1C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6792 0 0
2
5.89815e-315 5.53747e-315
0
14 Logic Display~
6 1270 2503 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L13
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
5.89815e-315 5.53812e-315
0
14 Logic Display~
6 1362 2512 0 1 2
10 34
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L14
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6316 0 0
2
5.89815e-315 5.53877e-315
0
9 Inverter~
13 1301 2375 0 2 22
0 54 25
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U4A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
8734 0 0
2
5.89815e-315 5.53941e-315
0
14 Logic Display~
6 1304 2514 0 1 2
10 25
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L15
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7988 0 0
2
5.89815e-315 5.54006e-315
0
14 Logic Display~
6 1409 2210 0 1 2
10 104
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L16
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3217 0 0
2
5.89815e-315 5.54071e-315
0
14 Logic Display~
6 1410 2185 0 1 2
10 103
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L17
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3965 0 0
2
5.89815e-315 5.54136e-315
0
14 Logic Display~
6 1407 2154 0 1 2
10 101
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L18
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8239 0 0
2
5.89815e-315 5.542e-315
0
14 Logic Display~
6 1411 2133 0 1 2
10 96
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L19
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
828 0 0
2
5.89815e-315 5.54265e-315
0
14 Logic Display~
6 1409 2104 0 1 2
10 94
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L20
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
5.89815e-315 5.5433e-315
0
14 Logic Display~
6 1407 2074 0 1 2
10 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L21
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7107 0 0
2
5.89815e-315 5.54395e-315
0
14 Logic Display~
6 1407 2044 0 1 2
10 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6433 0 0
2
5.89815e-315 5.54459e-315
0
14 Logic Display~
6 1409 2006 0 1 2
10 6
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L23
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8559 0 0
2
5.89815e-315 5.54524e-315
0
14 Logic Display~
6 1409 1970 0 1 2
10 100
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L24
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3674 0 0
2
5.89815e-315 5.54589e-315
0
14 Logic Display~
6 1235 1919 0 1 2
10 60
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L25
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5697 0 0
2
5.89815e-315 5.54654e-315
0
14 Logic Display~
6 1234 1889 0 1 2
10 88
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L26
40 4 61 12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
5.89815e-315 5.54719e-315
0
14 Logic Display~
6 1260 1871 0 1 2
10 9
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L27
-8 -21 13 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5219 0 0
2
5.89815e-315 5.54783e-315
0
14 Logic Display~
6 1234 1841 0 1 2
10 93
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L28
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3795 0 0
2
5.89815e-315 5.54848e-315
0
14 Logic Display~
6 1098 2498 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L35
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3637 0 0
2
5.89815e-315 5.54978e-315
0
5 4025~
219 621 2291 0 4 22
0 91 131 60 86
0
0 0 624 270
4 4025
-14 -24 14 -16
3 U2A
35 -10 56 -2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 512 3 1 2 0
1 U
3226 0 0
2
5.89815e-315 5.55042e-315
0
7 74LS126
116 600 269 0 12 25
0 60 110 60 109 60 108 60 107 30
31 32 33
0
0 0 4848 0
7 74LS126
-24 -51 25 -43
3 U17
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
6966 0 0
2
5.89815e-315 5.55107e-315
0
7 74LS193
137 429 266 0 14 29
0 88 89 87 2 30 31 32 33 132
133 110 109 108 107
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U16
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9796 0 0
2
5.89815e-315 5.55172e-315
0
14 Logic Display~
6 737 168 0 1 2
10 70
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L29
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
5.89815e-315 5.55237e-315
0
14 Logic Display~
6 769 168 0 1 2
10 69
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L30
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
5.89815e-315 5.55301e-315
0
14 Logic Display~
6 807 168 0 1 2
10 68
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L31
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
5.89815e-315 5.55366e-315
0
14 Logic Display~
6 846 166 0 1 2
10 67
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L32
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
5.89815e-315 5.55398e-315
0
14 Logic Display~
6 885 165 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L33
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4681 0 0
2
5.89815e-315 5.55431e-315
0
14 Logic Display~
6 922 165 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L34
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9730 0 0
2
5.89815e-315 5.55463e-315
0
14 Logic Display~
6 961 164 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L36
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9874 0 0
2
5.89815e-315 5.55496e-315
0
14 Logic Display~
6 1003 166 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L37
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
364 0 0
2
5.89815e-315 5.55528e-315
0
295
14 0 3 0 0 16512 0 35 0 0 219 6
1200 691
1175 691
1175 767
1624 767
1624 2381
1150 2381
2 0 4 0 0 8320 0 35 0 0 4 5
1264 691
1675 691
1675 2317
1414 2317
1414 2339
0 3 5 0 0 8320 0 0 35 5 0 4
1446 2329
1607 2329
1607 682
1264 682
0 1 4 0 0 0 0 0 16 263 0 5
1229 2078
1229 2339
1422 2339
1422 2523
1423 2523
3 1 5 0 0 0 0 17 15 0 0 4
1446 2315
1446 2499
1529 2499
1529 2518
1 0 3 0 0 0 0 17 0 0 264 4
1455 2269
1455 2241
1310 2241
1310 2048
2 0 4 0 0 0 0 17 0 0 263 3
1437 2269
1292 2269
1292 2078
1 0 6 0 0 4096 0 109 0 0 9 2
1270 2489
1270 2094
0 0 6 0 0 0 0 0 0 0 265 3
1280 2094
1244 2094
1244 2010
2 0 3 0 0 0 0 106 0 0 264 2
1188 2244
1188 2048
1 3 7 0 0 4224 0 18 19 0 0 3
366 1632
366 1645
361 1645
1 0 8 0 0 4096 0 1 0 0 204 2
308 1720
156 1720
2 0 9 0 0 4096 0 108 0 0 275 4
1320 2250
1320 1944
1066 1944
1066 1875
13 1 10 0 0 4224 0 67 80 0 0 3
253 1944
253 2214
327 2214
1 14 11 0 0 8320 0 79 67 0 0 3
326 2189
244 2189
244 1944
1 15 12 0 0 8320 0 78 67 0 0 3
328 2158
235 2158
235 1944
1 16 13 0 0 8320 0 77 67 0 0 3
328 2136
226 2136
226 1944
1 17 14 0 0 8320 0 76 67 0 0 3
328 2108
217 2108
217 1944
1 18 15 0 0 8320 0 75 67 0 0 3
330 2078
208 2078
208 1944
1 19 16 0 0 4224 0 74 67 0 0 3
332 2048
199 2048
199 1944
1 20 17 0 0 4224 0 73 67 0 0 3
332 2010
190 2010
190 1944
1 21 18 0 0 4224 0 72 67 0 0 3
332 1974
181 1974
181 1944
0 1 19 0 0 8320 0 0 23 83 0 4
1137 601
1137 546
1246 546
1246 520
0 1 20 0 0 8320 0 0 22 82 0 4
1169 610
1169 559
1277 559
1277 518
0 1 21 0 0 8320 0 0 21 81 0 4
1185 619
1185 529
1310 529
1310 516
0 1 22 0 0 8320 0 0 20 80 0 4
1178 628
1178 537
1342 537
1342 516
1 0 23 0 0 0 0 24 0 0 94 2
1529 430
1529 430
10 9 24 0 0 4096 0 30 30 0 0 2
1256 1406
1265 1406
9 0 24 0 0 4096 0 30 0 0 30 2
1265 1406
1329 1406
1 0 24 0 0 8320 0 30 0 0 0 3
1265 1336
1329 1336
1329 1417
2 0 25 0 0 4096 0 30 0 0 32 2
1256 1330
1256 1301
3 0 25 0 0 12416 0 30 0 0 213 5
1247 1330
1247 1301
1619 1301
1619 2484
1304 2484
4 0 8 0 0 8192 0 30 0 0 287 3
1238 1336
1238 1291
1724 1291
11 1 26 0 0 8320 0 30 28 0 0 4
1229 1400
1229 1494
1403 1494
1403 1396
12 1 27 0 0 8320 0 30 27 0 0 4
1220 1400
1220 1475
1431 1475
1431 1397
13 1 28 0 0 8320 0 30 26 0 0 4
1211 1400
1211 1463
1461 1463
1461 1396
14 1 29 0 0 8320 0 30 25 0 0 5
1202 1400
1202 1450
1483 1450
1483 1392
1484 1392
5 0 30 0 0 8192 0 30 0 0 291 3
1229 1336
1229 1290
885 1290
6 0 31 0 0 8192 0 30 0 0 290 3
1220 1336
1220 1308
922 1308
7 0 32 0 0 8192 0 30 0 0 289 3
1211 1336
1211 1325
961 1325
8 0 33 0 0 4096 0 30 0 0 288 2
1202 1336
1003 1336
1 0 34 0 0 4096 0 33 0 0 45 2
1092 959
1097 959
3 0 34 0 0 0 0 33 0 0 45 2
1092 941
1097 941
5 0 34 0 0 0 0 33 0 0 45 2
1092 923
1097 923
0 7 34 0 0 8320 0 0 33 214 0 6
1329 2359
1628 2359
1628 973
1097 973
1097 905
1092 905
2 0 35 0 0 4224 0 33 0 0 57 2
1092 950
1289 950
4 0 36 0 0 4224 0 33 0 0 56 2
1092 932
1307 932
6 0 37 0 0 4224 0 33 0 0 55 2
1092 914
1325 914
8 0 38 0 0 4224 0 33 0 0 54 2
1092 896
1343 896
9 1 39 0 0 8320 0 34 2 0 0 5
1352 871
1352 1043
1555 1043
1555 1101
1554 1101
7 1 40 0 0 8320 0 34 3 0 0 5
1334 871
1334 1024
1523 1024
1523 1101
1521 1101
5 1 41 0 0 8320 0 34 4 0 0 5
1316 871
1316 1003
1486 1003
1486 1101
1484 1101
3 1 42 0 0 8320 0 34 5 0 0 5
1298 871
1298 991
1451 991
1451 1099
1449 1099
8 1 38 0 0 0 0 34 6 0 0 5
1343 871
1343 1042
1229 1042
1229 1098
1228 1098
6 1 37 0 0 0 0 34 7 0 0 5
1325 871
1325 1023
1190 1023
1190 1096
1188 1096
4 1 36 0 0 0 0 34 8 0 0 5
1307 871
1307 1003
1152 1003
1152 1096
1150 1096
2 1 35 0 0 0 0 34 9 0 0 5
1289 871
1289 991
1114 991
1114 1095
1113 1095
2 1 43 0 0 12416 0 32 34 0 0 6
1378 2293
1378 2391
1639 2391
1639 889
1280 889
1280 871
0 1 3 0 0 0 0 0 32 264 0 2
1378 2048
1378 2257
10 1 2 0 0 4096 0 34 31 0 0 2
1361 877
1443 877
9 11 44 0 0 8320 0 35 34 0 0 3
1270 628
1298 628
1298 807
10 12 45 0 0 8320 0 35 34 0 0 3
1270 619
1316 619
1316 807
11 13 46 0 0 8320 0 35 34 0 0 3
1270 610
1334 610
1334 807
12 14 47 0 0 8320 0 35 34 0 0 3
1270 601
1352 601
1352 807
9 0 30 0 0 0 0 33 0 0 291 4
1028 950
900 950
900 945
885 945
10 0 31 0 0 0 0 33 0 0 290 4
1028 932
937 932
937 927
922 927
11 0 32 0 0 0 0 33 0 0 289 4
1028 914
976 914
976 909
961 909
12 0 33 0 0 0 0 33 0 0 288 4
1028 896
1014 896
1014 891
1003 891
13 0 6 0 0 16512 0 35 0 0 8 6
1200 700
1186 700
1186 743
1649 743
1649 2468
1270 2468
1 0 48 0 0 16512 0 35 0 0 217 6
1264 700
1604 700
1604 717
1662 717
1662 2397
1209 2397
4 0 6 0 0 8320 0 35 0 0 209 4
1264 673
1685 673
1685 2420
1098 2420
5 0 49 0 0 8192 0 35 0 0 95 3
1270 664
1419 664
1419 444
6 0 50 0 0 8320 0 35 0 0 96 3
1270 655
1409 655
1409 435
7 0 51 0 0 8192 0 35 0 0 97 3
1270 646
1401 646
1401 426
8 0 52 0 0 8320 0 35 0 0 98 3
1270 637
1392 637
1392 417
3 0 53 0 0 4096 0 36 0 0 79 2
1123 643
1153 643
5 0 53 0 0 0 0 36 0 0 79 2
1123 625
1153 625
7 0 53 0 0 0 0 36 0 0 79 2
1123 607
1153 607
1 0 53 0 0 16512 0 36 0 0 220 6
1123 661
1153 661
1153 572
1694 572
1694 2429
1047 2429
2 19 22 0 0 0 0 36 35 0 0 4
1123 652
1169 652
1169 628
1194 628
4 20 21 0 0 0 0 36 35 0 0 4
1123 634
1166 634
1166 619
1194 619
6 21 20 0 0 0 0 36 35 0 0 4
1123 616
1159 616
1159 610
1194 610
8 22 19 0 0 0 0 36 35 0 0 3
1123 598
1123 601
1194 601
9 0 30 0 0 0 0 36 0 0 291 2
1059 652
885 652
10 0 31 0 0 0 0 36 0 0 290 2
1059 634
922 634
11 0 32 0 0 0 0 36 0 0 289 2
1059 616
961 616
12 0 33 0 0 0 0 36 0 0 288 2
1059 598
1003 598
0 1 52 0 0 0 0 0 37 110 0 3
1130 368
1321 368
1321 212
0 1 51 0 0 4224 0 0 38 109 0 3
1139 358
1371 358
1371 218
0 1 50 0 0 0 0 0 39 108 0 4
1148 352
1339 352
1339 221
1416 221
0 1 49 0 0 4224 0 0 40 107 0 3
1157 344
1438 344
1438 220
9 0 2 0 0 0 0 44 0 0 93 3
1193 338
1262 338
1262 302
1 1 2 0 0 0 0 44 42 0 0 4
1193 268
1253 268
1253 302
1275 302
5 1 23 0 0 28800 0 41 83 0 0 9
1500 430
1569 430
1569 1016
1589 1016
1589 1124
1549 1124
1549 1816
520 1816
520 2227
0 4 49 0 0 0 0 0 41 107 0 4
1157 425
1291 425
1291 444
1444 444
0 3 50 0 0 0 0 0 41 108 0 4
1148 409
1305 409
1305 435
1444 435
0 2 51 0 0 0 0 0 41 109 0 4
1139 385
1318 385
1318 426
1444 426
0 1 52 0 0 0 0 0 41 110 0 4
1130 380
1331 380
1331 417
1444 417
9 0 30 0 0 0 0 43 0 0 291 2
1047 440
885 440
10 0 31 0 0 0 0 43 0 0 290 2
1047 422
922 422
11 0 32 0 0 0 0 43 0 0 289 2
1047 404
961 404
12 0 33 0 0 0 0 43 0 0 288 2
1047 386
1003 386
1 0 54 0 0 4096 0 43 0 0 106 3
1111 449
1170 449
1170 395
3 0 54 0 0 0 0 43 0 0 106 3
1111 431
1143 431
1143 395
5 0 54 0 0 0 0 43 0 0 106 3
1111 413
1129 413
1129 395
7 0 54 0 0 8320 0 43 0 0 226 4
1111 395
1702 395
1702 2441
980 2441
2 11 49 0 0 0 0 43 44 0 0 3
1111 440
1157 440
1157 332
4 12 50 0 0 0 0 43 44 0 0 3
1111 422
1148 422
1148 332
6 13 51 0 0 0 0 43 44 0 0 3
1111 404
1139 404
1139 332
8 14 52 0 0 0 0 43 44 0 0 3
1111 386
1130 386
1130 332
2 0 55 0 0 4096 0 44 0 0 112 2
1184 262
1184 227
3 0 55 0 0 12416 0 44 0 0 229 5
1175 262
1175 227
1712 227
1712 2453
895 2453
10 9 2 0 0 0 0 44 44 0 0 2
1184 338
1193 338
4 0 8 0 0 0 0 44 0 0 287 2
1166 268
1166 59
5 0 30 0 0 0 0 44 0 0 291 3
1157 268
1157 228
885 228
6 0 31 0 0 0 0 44 0 0 290 3
1148 268
1148 240
922 240
7 0 32 0 0 0 0 44 0 0 289 3
1139 268
1139 255
961 255
8 0 33 0 0 0 0 44 0 0 288 2
1130 268
1003 268
14 3 56 0 0 12416 0 58 67 0 0 4
303 1326
303 1449
226 1449
226 1874
4 13 57 0 0 4224 0 67 58 0 0 4
217 1874
217 1437
312 1437
312 1326
5 12 58 0 0 4224 0 67 58 0 0 4
208 1874
208 1418
321 1418
321 1326
6 11 59 0 0 4224 0 67 58 0 0 4
199 1874
199 1401
330 1401
330 1326
1 1 2 0 0 0 0 53 54 0 0 2
457 1660
457 1661
2 0 60 0 0 8192 0 54 0 0 277 3
475 1661
651 1661
651 1923
1 3 61 0 0 12416 0 58 54 0 0 4
366 1262
366 1257
466 1257
466 1612
12 0 30 0 0 0 0 56 0 0 291 2
694 1485
885 1485
11 0 31 0 0 0 0 56 0 0 290 2
694 1467
922 1467
10 0 32 0 0 4096 0 56 0 0 289 2
694 1449
961 1449
9 0 33 0 0 4096 0 56 0 0 288 2
694 1431
1003 1431
5 0 62 0 0 4096 0 56 0 0 133 2
630 1458
566 1458
3 0 62 0 0 0 0 56 0 0 133 2
630 1440
566 1440
1 0 62 0 0 0 0 56 0 0 133 2
630 1422
566 1422
7 0 62 0 0 16512 0 56 0 0 238 6
630 1476
566 1476
566 1387
79 1387
79 2444
836 2444
14 8 63 0 0 4224 0 57 56 0 0 3
510 1326
510 1485
630 1485
13 6 64 0 0 4224 0 57 56 0 0 3
519 1326
519 1467
630 1467
12 4 65 0 0 4224 0 57 56 0 0 3
528 1326
528 1449
630 1449
11 2 66 0 0 4224 0 57 56 0 0 3
537 1326
537 1431
630 1431
5 0 33 0 0 8192 0 57 0 0 288 3
537 1262
537 1233
1003 1233
6 0 32 0 0 8192 0 57 0 0 289 3
528 1262
528 1214
961 1214
7 0 31 0 0 8192 0 57 0 0 290 3
519 1262
519 1203
922 1203
8 0 30 0 0 8192 0 57 0 0 291 3
510 1262
510 1189
885 1189
5 0 67 0 0 8192 0 58 0 0 292 3
330 1262
330 1179
846 1179
6 0 68 0 0 8192 0 58 0 0 293 3
321 1262
321 1166
807 1166
7 0 69 0 0 8192 0 58 0 0 294 3
312 1262
312 1149
769 1149
0 0 70 0 0 8192 0 0 0 0 295 3
302 1268
302 1127
737 1127
3 0 71 0 0 4096 0 58 0 0 149 2
348 1256
348 1219
2 0 71 0 0 0 0 58 0 0 149 2
357 1256
357 1219
3 0 71 0 0 0 0 57 0 0 149 2
555 1256
555 1219
2 0 71 0 0 12416 0 57 0 0 241 5
564 1256
564 1219
96 1219
96 2426
786 2426
10 0 2 0 0 0 0 58 0 0 151 3
357 1332
357 1338
366 1338
9 0 2 0 0 8320 0 58 0 0 154 4
366 1332
366 1339
628 1339
628 1332
10 9 2 0 0 0 0 57 57 0 0 2
564 1332
573 1332
0 1 2 0 0 0 0 0 55 154 0 2
663 1332
663 1342
9 0 2 0 0 0 0 57 0 0 155 2
573 1332
663 1332
1 0 2 0 0 0 0 57 0 0 0 4
573 1262
573 1241
663 1241
663 1337
0 4 8 0 0 0 0 0 57 157 0 3
339 1194
546 1194
546 1262
4 0 8 0 0 0 0 58 0 0 204 3
339 1262
339 1194
156 1194
1 0 72 0 0 8320 0 60 0 0 243 4
564 917
106 917
106 2386
721 2386
14 0 33 0 0 0 0 60 0 0 288 2
634 989
1003 989
13 0 32 0 0 0 0 60 0 0 289 2
634 980
961 980
12 0 31 0 0 0 0 60 0 0 290 2
634 971
922 971
11 0 30 0 0 0 0 60 0 0 291 2
634 962
885 962
10 0 67 0 0 0 0 60 0 0 292 2
634 953
846 953
9 0 68 0 0 0 0 60 0 0 293 2
634 944
807 944
8 0 69 0 0 0 0 60 0 0 294 2
634 935
769 935
7 0 70 0 0 0 0 60 0 0 295 2
634 926
737 926
2 1 2 0 0 0 0 60 59 0 0 2
570 953
372 953
14 3 73 0 0 8320 0 63 60 0 0 3
420 834
420 962
570 962
13 4 74 0 0 4224 0 63 60 0 0 3
438 834
438 971
570 971
12 5 75 0 0 4224 0 63 60 0 0 3
456 834
456 980
570 980
11 6 76 0 0 4224 0 63 60 0 0 3
474 834
474 989
570 989
10 1 2 0 0 0 0 63 61 0 0 4
411 764
411 734
378 734
378 736
9 1 77 0 0 8320 0 63 13 0 0 5
420 770
420 634
209 634
209 688
200 688
3 1 78 0 0 8320 0 63 10 0 0 5
474 770
474 688
291 688
291 766
276 766
5 1 79 0 0 8320 0 63 11 0 0 5
456 770
456 667
258 667
258 745
245 745
7 1 80 0 0 8320 0 63 12 0 0 5
438 770
438 648
227 648
227 724
213 724
1 1 81 0 0 8320 0 63 14 0 0 5
492 770
492 619
214 619
214 600
213 600
2 11 82 0 0 4224 0 63 64 0 0 4
483 770
483 648
564 648
564 631
12 4 83 0 0 12416 0 64 63 0 0 4
555 631
555 642
465 642
465 770
6 13 84 0 0 4224 0 63 64 0 0 4
447 770
447 636
546 636
546 631
14 8 85 0 0 8320 0 64 63 0 0 3
537 631
429 631
429 770
10 0 2 0 0 0 0 64 0 0 184 4
591 637
591 647
656 647
656 567
9 0 2 0 0 0 0 64 0 0 184 3
600 637
669 637
669 567
1 1 2 0 0 0 0 64 62 0 0 4
600 567
681 567
681 587
685 587
2 0 86 0 0 4096 0 64 0 0 186 3
591 561
591 496
582 496
3 0 86 0 0 12416 0 64 0 0 248 5
582 561
582 484
143 484
143 2367
627 2367
4 0 8 0 0 0 0 64 0 0 204 3
573 567
573 497
156 497
5 0 33 0 0 0 0 64 0 0 288 3
564 567
564 557
1003 557
6 0 32 0 0 0 0 64 0 0 289 3
555 567
555 547
961 547
7 0 31 0 0 0 0 64 0 0 290 3
546 567
546 531
922 531
8 0 30 0 0 0 0 64 0 0 291 3
537 567
537 517
885 517
8 0 33 0 0 12288 0 129 0 0 288 4
397 302
378 302
378 363
1003 363
7 0 32 0 0 12288 0 129 0 0 289 4
397 293
364 293
364 346
961 346
6 0 31 0 0 12288 0 129 0 0 290 4
397 284
351 284
351 333
922 333
5 0 30 0 0 12288 0 129 0 0 291 4
397 275
338 275
338 321
885 321
0 3 87 0 0 8320 0 0 129 252 0 4
493 2432
126 2432
126 257
391 257
1 0 88 0 0 8320 0 129 0 0 257 4
397 239
138 239
138 2230
425 2230
4 1 2 0 0 0 0 129 65 0 0 3
397 266
339 266
339 180
2 1 89 0 0 8320 0 129 66 0 0 3
397 248
364 248
364 178
5 0 60 0 0 0 0 128 0 0 203 2
568 278
548 278
3 0 60 0 0 0 0 128 0 0 203 2
568 260
548 260
1 0 60 0 0 0 0 128 0 0 203 2
568 242
548 242
0 7 60 0 0 8320 0 0 128 208 0 6
387 2401
117 2401
117 200
548 200
548 296
568 296
3 0 8 0 0 16512 0 68 0 0 287 5
380 1860
331 1860
331 1846
156 1846
156 59
3 1 90 0 0 8320 0 84 85 0 0 4
500 2336
504 2336
504 2374
502 2374
1 3 91 0 0 4224 0 127 87 0 0 2
636 2272
636 2273
0 0 60 0 0 0 0 0 0 277 208 6
478 1923
478 1940
378 1940
378 2377
387 2377
387 2393
0 1 60 0 0 0 0 0 81 0 0 2
387 2388
387 2465
0 1 6 0 0 0 0 0 126 225 0 5
1064 2029
1089 2029
1089 2399
1098 2399
1098 2484
0 0 92 0 0 4224 0 0 0 0 0 3
511 2460
511 2461
512 2461
1 0 93 0 0 4096 0 125 0 0 274 2
1218 1845
1218 1868
1 0 88 0 0 0 0 123 0 0 276 2
1218 1893
1218 1893
2 1 25 0 0 0 0 111 112 0 0 2
1304 2393
1304 2500
3 1 34 0 0 0 0 108 110 0 0 3
1329 2295
1329 2498
1362 2498
0 1 54 0 0 0 0 0 111 226 0 3
980 2360
1304 2360
1304 2357
1 0 94 0 0 4096 0 108 0 0 262 2
1338 2250
1338 2108
3 1 48 0 0 0 0 106 107 0 0 6
1197 2290
1197 2321
1188 2321
1188 2349
1209 2349
1209 2483
1 0 6 0 0 0 0 106 0 0 265 2
1206 2244
1206 2010
0 1 3 0 0 0 0 0 105 264 0 4
1130 2048
1130 2301
1150 2301
1150 2467
3 1 53 0 0 0 0 103 104 0 0 2
1047 2353
1047 2477
4 1 95 0 0 8320 0 102 103 0 0 3
1055 2288
1056 2288
1056 2308
0 2 9 0 0 0 0 0 103 227 0 3
971 2225
1038 2225
1038 2308
3 0 4 0 0 0 0 102 0 0 263 2
1046 2242
1046 2078
2 0 3 0 0 0 0 102 0 0 264 2
1055 2243
1055 2048
1 0 6 0 0 0 0 102 0 0 265 2
1064 2242
1064 2010
3 1 54 0 0 0 0 100 101 0 0 2
980 2283
980 2467
0 2 9 0 0 0 0 0 100 232 0 3
890 2044
971 2044
971 2238
1 0 96 0 0 4096 0 100 0 0 261 2
989 2238
989 2136
1 3 55 0 0 0 0 99 98 0 0 4
895 2475
895 2416
896 2416
896 2417
0 2 97 0 0 12416 0 0 98 247 0 5
730 2293
795 2293
795 2339
887 2339
887 2365
3 1 98 0 0 4224 0 97 98 0 0 3
899 2341
899 2365
905 2365
0 2 9 0 0 0 0 0 97 239 0 3
809 2036
890 2036
890 2296
1 5 99 0 0 4224 0 97 96 0 0 2
908 2296
908 2284
4 0 94 0 0 0 0 96 0 0 262 2
894 2234
894 2108
3 0 4 0 0 0 0 96 0 0 263 2
903 2234
903 2078
2 0 3 0 0 0 0 96 0 0 264 2
912 2234
912 2048
1 0 6 0 0 0 0 96 0 0 265 2
921 2234
921 2010
3 1 62 0 0 0 0 94 95 0 0 4
818 2328
818 2343
836 2343
836 2470
0 2 9 0 0 0 0 0 94 250 0 3
627 2020
809 2020
809 2277
0 1 100 0 0 8192 0 0 94 246 0 5
739 2002
818 2002
818 2271
827 2271
827 2277
1 2 71 0 0 0 0 93 92 0 0 4
786 2467
786 2389
787 2389
787 2390
0 0 88 0 0 0 0 0 0 257 0 2
425 2355
787 2355
3 1 72 0 0 0 0 89 91 0 0 2
721 2351
721 2467
0 2 88 0 0 0 0 0 89 257 0 3
425 2147
712 2147
712 2299
2 0 93 0 0 4096 0 88 0 0 274 2
721 2232
721 1868
0 1 100 0 0 0 0 0 88 251 0 3
645 1991
739 1991
739 2232
1 3 97 0 0 0 0 89 88 0 0 2
730 2299
730 2277
4 1 86 0 0 0 0 127 90 0 0 2
627 2324
627 2474
3 0 60 0 0 0 0 127 0 0 277 2
618 2272
618 1923
0 2 9 0 0 0 0 0 87 253 0 3
482 1964
627 1964
627 2228
1 0 100 0 0 0 0 87 0 0 266 2
645 2228
645 1974
3 1 87 0 0 0 0 85 86 0 0 2
493 2425
493 2458
2 0 9 0 0 4096 0 85 0 0 275 6
484 2374
484 1964
482 1964
482 1949
516 1949
516 1878
1 0 101 0 0 4096 0 84 0 0 260 2
491 2290
491 2158
2 3 102 0 0 8320 0 84 83 0 0 5
509 2290
522 2290
522 2266
511 2266
511 2272
2 0 103 0 0 4096 0 83 0 0 259 4
502 2227
502 2204
500 2204
500 2189
0 1 88 0 0 0 0 0 82 276 0 6
494 1893
494 1908
425 1908
425 2355
428 2355
428 2480
2 1 104 0 0 4224 0 80 113 0 0 2
363 2214
1393 2214
2 1 103 0 0 4224 0 79 114 0 0 2
362 2189
1394 2189
2 1 101 0 0 4224 0 78 115 0 0 2
364 2158
1391 2158
2 1 96 0 0 4224 0 77 116 0 0 3
364 2136
1395 2136
1395 2137
2 1 94 0 0 4224 0 76 117 0 0 2
364 2108
1393 2108
2 1 4 0 0 128 0 75 118 0 0 2
366 2078
1391 2078
2 1 3 0 0 0 0 74 119 0 0 2
368 2048
1391 2048
2 1 6 0 0 0 0 73 120 0 0 2
368 2010
1393 2010
2 1 100 0 0 4224 0 72 121 0 0 2
368 1974
1393 1974
1 0 2 0 0 0 0 67 0 0 268 2
262 1868
262 1861
1 2 2 0 0 0 0 71 67 0 0 3
287 1861
253 1861
253 1868
3 0 9 0 0 0 0 70 0 0 275 5
304 1834
280 1834
280 1785
480 1785
480 1878
2 0 88 0 0 0 0 70 0 0 276 5
305 1825
286 1825
286 1790
470 1790
470 1893
1 0 60 0 0 0 0 70 0 0 277 5
304 1816
292 1816
292 1794
461 1794
461 1923
0 2 105 0 0 4224 0 0 68 273 0 3
370 1823
370 1842
380 1842
4 1 105 0 0 0 0 70 68 0 0 6
356 1825
370 1825
370 1823
382 1823
382 1833
380 1833
9 0 93 0 0 8320 0 68 0 0 0 3
444 1869
444 1868
1222 1868
10 1 9 0 0 12416 0 68 124 0 0 4
444 1878
516 1878
516 1875
1244 1875
11 0 88 0 0 0 0 68 0 0 0 3
444 1887
444 1893
1222 1893
12 1 60 0 0 0 0 68 122 0 0 3
444 1896
444 1923
1219 1923
1 4 106 0 0 4224 0 69 68 0 0 4
359 1881
370 1881
370 1878
374 1878
12 0 33 0 0 0 0 128 0 0 288 2
632 305
1003 305
11 0 32 0 0 0 0 128 0 0 289 2
632 287
961 287
10 0 31 0 0 0 0 128 0 0 290 2
632 269
922 269
9 0 30 0 0 0 0 128 0 0 291 2
632 251
885 251
14 8 107 0 0 8320 0 129 128 0 0 3
461 302
461 305
568 305
13 6 108 0 0 4224 0 129 128 0 0 4
461 293
524 293
524 287
568 287
12 4 109 0 0 12416 0 129 128 0 0 4
461 284
507 284
507 269
568 269
11 2 110 0 0 12416 0 129 128 0 0 4
461 275
488 275
488 251
568 251
0 0 8 0 0 0 0 0 0 0 0 3
124 59
1724 59
1724 1583
1 1 33 0 0 4224 0 137 45 0 0 3
1003 184
1003 1657
1004 1657
1 1 32 0 0 4224 0 136 46 0 0 2
961 182
961 1654
1 1 31 0 0 4224 0 135 47 0 0 2
922 183
922 1651
1 1 30 0 0 4224 0 134 48 0 0 3
885 183
885 1649
886 1649
1 1 67 0 0 4224 0 133 49 0 0 2
846 184
846 1650
1 1 68 0 0 4224 0 132 50 0 0 2
807 186
807 1649
1 1 69 0 0 4224 0 131 51 0 0 2
769 186
769 1648
1 1 70 0 0 4224 0 130 52 0 0 2
737 186
737 1656
65
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
126 17 186 49
139 26 172 48
3 clk
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
279 1948 333 1980
289 1956 322 1978
3 LDA
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
282 1981 336 2013
292 1989 325 2011
3 ADD
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
283 2020 337 2052
293 2028 326 2050
3 SUB
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
282 2050 336 2082
292 2058 325 2080
3 AND
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
279 2076 333 2108
289 2084 322 2106
3 MOV
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
278 2103 332 2135
288 2111 321 2133
3 OUT
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
279 2128 333 2160
289 2136 322 2158
3 JMP
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
283 2161 326 2193
293 2169 315 2191
2 JZ
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
279 2186 333 2218
289 2194 322 2216
3 HLT
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
847 1917 890 1949
857 1925 879 1947
2 T1
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
794 1887 837 1919
804 1895 826 1917
2 T2
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
793 1836 836 1868
803 1844 825 1866
2 T4
-19 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
356 2485 406 2519
366 2493 395 2517
2 Ep
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
408 2498 459 2532
418 2506 448 2530
2 Cp
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
473 2489 524 2523
483 2497 513 2521
2 Lp
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
597 2497 654 2531
607 2505 643 2529
2 Lm
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
695 2508 750 2542
705 2516 739 2540
2 CE
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
760 2508 805 2542
770 2516 794 2540
2 Li
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
879 2506 929 2540
889 2514 918 2538
2 La
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
951 2506 1002 2540
961 2514 991 2538
2 Ea
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1028 2509 1080 2543
1038 2517 1069 2541
2 Eu
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1192 2519 1242 2553
1202 2527 1231 2551
2 S3
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1419 2550 1470 2584
1429 2558 1459 2582
2 S2
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1501 2551 1548 2585
1511 2559 1537 2583
2 S1
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1082 2521 1133 2555
1092 2529 1122 2553
2 S0
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
1233 2526 1294 2560
1244 2535 1282 2559
3 Cin
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1285 2523 1337 2557
1296 2532 1325 2556
2 Lo
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1348 2531 1402 2565
1359 2539 1390 2563
2 Eb
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
812 2503 861 2537
823 2511 849 2535
2 Ei
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
847 1868 888 1900
856 1877 878 1899
2 T3
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
228 163 277 195
241 171 263 193
2 Ep
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
229 211 278 243
242 220 264 242
2 Cp
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
230 251 279 283
243 259 265 281
2 Lp
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
478 131 553 179
492 140 538 174
2 PC
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 11
382 396 592 444
397 405 576 439
11 input & mar
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
254 446 305 478
268 454 290 476
2 Lm
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
178 536 306 568
192 545 291 567
9 SM(mar=1)
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
200 787 283 846
213 796 269 840
13 input 
SM=0
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
549 836 661 884
564 845 645 879
3 ROM
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
313 880 364 912
327 889 349 911
2 Cs
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
401 1054 473 1102
416 1063 457 1097
2 IR
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
400 1223 449 1255
413 1232 435 1254
2 Li
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
188 1352 237 1384
201 1361 223 1383
2 Ei
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 14
753 1765 992 1813
768 1774 976 1808
14 control matrix
-19 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1138 2501 1178 2535
1147 2510 1168 2534
1 M
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1469 195 1508 229
1477 201 1499 223
2 La
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1401 365 1440 399
1409 370 1431 392
2 Ea
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1225 112 1265 163
1234 117 1255 152
1 A
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1623 22 1683 54
1636 31 1669 53
3 clk
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
1106 494 1186 545
1112 499 1179 534
3 ALU
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1418 533 1457 567
1426 539 1448 561
2 Eu
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1495 440 1523 474
1503 445 1514 467
1 z
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1438 645 1477 679
1446 650 1468 672
2 S0
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1427 579 1466 613
1435 585 1457 607
2 S1
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1619 689 1658 723
1627 694 1649 716
2 S2
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1128 692 1156 726
1136 697 1147 719
1 M
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1447 698 1486 732
1455 704 1477 726
2 S3
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1364 743 1414 777
1372 748 1405 770
3 Cin
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1619 859 1647 893
1627 864 1638 886
1 S
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1105 1126 1149 1177
1114 1131 1139 1166
1 B
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1439 1130 1480 1181
1448 1135 1470 1170
1 C
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1363 945 1398 979
1369 950 1391 972
2 Eb
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 6
1269 1211 1380 1262
1278 1217 1370 1252
6 output
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1482 1296 1521 1330
1490 1302 1512 1324
2 Lo
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
