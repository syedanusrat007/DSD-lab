CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
48
13 Logic Switch~
5 145 315 0 1 11
0 23
0
0 0 21360 0
2 0V
-7 -16 7 -8
3 V48
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7479 0 0
2
42919.8 28
0
13 Logic Switch~
5 166 324 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V47
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5690 0 0
2
42919.8 27
0
13 Logic Switch~
5 188 333 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V46
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5617 0 0
2
42919.8 26
0
13 Logic Switch~
5 207 342 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V45
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3903 0 0
2
42919.8 25
0
13 Logic Switch~
5 225 351 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V44
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4452 0 0
2
42919.8 24
0
13 Logic Switch~
5 238 360 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V43
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6282 0 0
2
42919.8 23
0
13 Logic Switch~
5 249 369 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V42
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7187 0 0
2
42919.8 22
0
13 Logic Switch~
5 254 378 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V41
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6866 0 0
2
42919.8 21
0
13 Logic Switch~
5 254 502 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V32
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7670 0 0
2
42919.8 8
0
13 Logic Switch~
5 249 493 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V31
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
951 0 0
2
42919.8 7
0
13 Logic Switch~
5 238 484 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V30
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9536 0 0
2
42919.8 6
0
13 Logic Switch~
5 225 475 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V29
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5495 0 0
2
42919.8 5
0
13 Logic Switch~
5 207 466 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V28
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8152 0 0
2
42919.8 4
0
13 Logic Switch~
5 188 457 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V27
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6223 0 0
2
42919.8 3
0
13 Logic Switch~
5 166 448 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V26
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5441 0 0
2
42919.8 2
0
13 Logic Switch~
5 145 439 0 1 11
0 16
0
0 0 21360 0
2 0V
-7 -16 7 -8
3 V25
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3189 0 0
2
42919.8 1
0
13 Logic Switch~
5 146 194 0 1 11
0 30
0
0 0 21360 0
2 0V
-7 -16 7 -8
3 V24
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8460 0 0
2
42919.8 13
0
13 Logic Switch~
5 167 203 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V23
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5179 0 0
2
42919.8 12
0
13 Logic Switch~
5 189 212 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V22
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3593 0 0
2
42919.8 11
0
13 Logic Switch~
5 208 221 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V21
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3928 0 0
2
42919.8 10
0
13 Logic Switch~
5 226 230 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
363 0 0
2
42919.8 9
0
13 Logic Switch~
5 239 239 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8132 0 0
2
42919.8 8
0
13 Logic Switch~
5 250 248 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
65 0 0
2
42919.8 7
0
13 Logic Switch~
5 255 257 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6609 0 0
2
42919.8 6
0
13 Logic Switch~
5 603 70 0 1 11
0 9
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8995 0 0
2
42919.8 0
0
13 Logic Switch~
5 481 97 0 1 11
0 6
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3918 0 0
2
42919.8 0
0
13 Logic Switch~
5 504 88 0 1 11
0 7
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7519 0 0
2
42919.8 0
0
13 Logic Switch~
5 528 79 0 1 11
0 8
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
377 0 0
2
42919.8 0
0
13 Logic Switch~
5 255 133 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8816 0 0
2
42919.8 0
0
13 Logic Switch~
5 250 124 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3877 0 0
2
42919.8 0
0
13 Logic Switch~
5 239 115 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
926 0 0
2
42919.8 0
0
13 Logic Switch~
5 226 106 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7262 0 0
2
42919.8 0
0
13 Logic Switch~
5 208 97 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5267 0 0
2
42919.8 0
0
13 Logic Switch~
5 189 88 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8838 0 0
2
42919.8 0
0
13 Logic Switch~
5 167 79 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7159 0 0
2
42919.8 0
0
13 Logic Switch~
5 146 70 0 1 11
0 38
0
0 0 21360 0
2 0V
-7 -16 7 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5812 0 0
2
42919.8 0
0
7 74LS151
20 301 342 0 14 29
0 23 22 21 20 19 3 2 2 9
8 7 6 18 17
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
331 0 0
2
42919.8 29
0
14 Logic Display~
6 560 365 0 1 2
10 18
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9604 0 0
2
42919.8 16
0
14 Logic Display~
6 560 393 0 1 2
10 17
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7518 0 0
2
42919.8 15
0
14 Logic Display~
6 560 517 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4832 0 0
2
42919.8 14
0
14 Logic Display~
6 560 489 0 1 2
10 11
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6798 0 0
2
42919.8 13
0
7 74LS151
20 301 466 0 14 29
0 16 15 14 13 12 2 5 5 9
8 7 6 11 10
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
3336 0 0
2
42919.8 0
0
7 74LS151
20 302 221 0 14 29
0 30 29 28 27 26 4 3 3 9
8 7 6 25 24
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
8370 0 0
2
42919.8 14
0
14 Logic Display~
6 561 244 0 1 2
10 25
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3910 0 0
2
42919.8 1
0
14 Logic Display~
6 561 272 0 1 2
10 24
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
316 0 0
2
42919.8 0
0
14 Logic Display~
6 561 148 0 1 2
10 31
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
536 0 0
2
42919.8 0
0
14 Logic Display~
6 561 120 0 1 2
10 32
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4460 0 0
2
42919.8 0
0
7 74LS151
20 302 97 0 14 29
0 38 37 36 35 34 33 4 4 9
8 7 6 32 31
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
3260 0 0
2
42919.8 0
0
118
8 6 2 0 0 4224 0 37 42 0 0 2
269 378
269 484
8 6 3 0 0 8320 0 43 37 0 0 3
270 257
269 257
269 360
8 6 4 0 0 4224 0 48 43 0 0 2
270 133
270 239
8 7 5 0 0 4096 0 42 42 0 0 2
269 502
269 493
8 7 2 0 0 0 0 37 37 0 0 2
269 378
269 369
8 7 3 0 0 0 0 43 43 0 0 2
270 257
270 248
8 7 4 0 0 0 0 48 48 0 0 2
270 133
270 124
0 0 6 0 0 4224 0 0 0 98 23 2
461 97
461 466
0 0 6 0 0 0 0 0 0 98 47 2
452 97
452 342
0 0 6 0 0 0 0 0 0 98 71 2
445 97
445 221
0 0 7 0 0 4224 0 0 0 99 24 2
439 88
439 457
0 0 7 0 0 0 0 0 0 99 48 2
427 88
427 333
0 0 7 0 0 0 0 0 0 99 72 2
416 88
416 212
0 0 8 0 0 4096 0 0 0 49 100 2
387 324
387 79
0 0 8 0 0 0 0 0 0 73 100 2
395 203
395 79
0 0 8 0 0 4224 0 0 0 25 100 2
408 448
408 79
0 0 9 0 0 4224 0 0 0 92 20 2
378 70
378 439
0 0 9 0 0 0 0 0 0 92 44 2
362 70
362 315
0 0 9 0 0 0 0 0 0 92 68 2
351 70
351 194
9 0 9 0 0 0 0 42 0 0 0 2
339 439
590 439
1 0 10 0 0 4096 0 40 0 0 26 2
544 521
544 502
1 0 11 0 0 0 0 41 0 0 27 2
544 493
544 493
12 0 6 0 0 0 0 42 0 0 0 2
333 466
488 466
11 0 7 0 0 0 0 42 0 0 0 2
333 457
510 457
10 0 8 0 0 0 0 42 0 0 0 2
333 448
531 448
14 0 10 0 0 4224 0 42 0 0 0 2
339 502
550 502
13 0 11 0 0 4224 0 42 0 0 0 2
333 493
549 493
1 0 5 0 0 0 0 9 0 0 36 2
266 502
266 502
1 0 5 0 0 0 0 10 0 0 37 2
261 493
261 493
1 0 2 0 0 0 0 11 0 0 38 2
250 484
250 484
1 0 12 0 0 0 0 12 0 0 39 2
237 475
237 475
1 0 13 0 0 0 0 13 0 0 40 2
219 466
219 466
1 0 14 0 0 0 0 14 0 0 41 2
200 457
200 457
1 0 15 0 0 0 0 15 0 0 42 2
178 448
178 448
1 0 16 0 0 0 0 16 0 0 43 2
157 439
157 439
8 0 5 0 0 4224 0 42 0 0 0 2
269 502
257 502
7 0 5 0 0 4224 0 42 0 0 0 2
269 493
249 493
6 0 2 0 0 128 0 42 0 0 0 2
269 484
235 484
5 0 12 0 0 4224 0 42 0 0 0 2
269 475
222 475
4 0 13 0 0 4224 0 42 0 0 0 2
269 466
204 466
3 0 14 0 0 4224 0 42 0 0 0 2
269 457
182 457
2 0 15 0 0 4224 0 42 0 0 0 2
269 448
160 448
1 0 16 0 0 4224 0 42 0 0 0 2
269 439
143 439
9 0 9 0 0 0 0 37 0 0 0 2
339 315
590 315
1 0 17 0 0 4096 0 39 0 0 50 2
544 397
544 378
1 0 18 0 0 0 0 38 0 0 51 2
544 369
544 369
12 0 6 0 0 0 0 37 0 0 0 2
333 342
488 342
11 0 7 0 0 0 0 37 0 0 0 2
333 333
510 333
10 0 8 0 0 0 0 37 0 0 0 2
333 324
531 324
14 0 17 0 0 4224 0 37 0 0 0 2
339 378
550 378
13 0 18 0 0 4224 0 37 0 0 0 2
333 369
549 369
1 0 2 0 0 0 0 8 0 0 60 2
266 378
266 378
1 0 2 0 0 0 0 7 0 0 61 2
261 369
261 369
1 0 3 0 0 0 0 6 0 0 62 2
250 360
250 360
1 0 19 0 0 0 0 5 0 0 63 2
237 351
237 351
1 0 20 0 0 0 0 4 0 0 64 2
219 342
219 342
1 0 21 0 0 0 0 3 0 0 65 2
200 333
200 333
1 0 22 0 0 0 0 2 0 0 66 2
178 324
178 324
1 0 23 0 0 0 0 1 0 0 67 2
157 315
157 315
8 0 2 0 0 144 0 37 0 0 5 2
269 378
257 378
7 0 2 0 0 128 0 37 0 0 5 2
269 369
249 369
6 0 3 0 0 128 0 37 0 0 0 2
269 360
235 360
5 0 19 0 0 4224 0 37 0 0 0 2
269 351
222 351
4 0 20 0 0 4224 0 37 0 0 0 2
269 342
204 342
3 0 21 0 0 4224 0 37 0 0 0 2
269 333
182 333
2 0 22 0 0 4224 0 37 0 0 0 2
269 324
160 324
1 0 23 0 0 4224 0 37 0 0 0 2
269 315
143 315
9 0 9 0 0 0 0 43 0 0 0 2
340 194
591 194
1 0 24 0 0 4096 0 45 0 0 74 2
545 276
545 257
1 0 25 0 0 0 0 44 0 0 75 2
545 248
545 248
12 0 6 0 0 0 0 43 0 0 0 2
334 221
489 221
11 0 7 0 0 0 0 43 0 0 0 2
334 212
511 212
10 0 8 0 0 0 0 43 0 0 0 2
334 203
532 203
14 0 24 0 0 4224 0 43 0 0 0 2
340 257
551 257
13 0 25 0 0 4224 0 43 0 0 0 2
334 248
550 248
1 0 3 0 0 0 0 24 0 0 84 2
267 257
267 257
1 0 3 0 0 0 0 23 0 0 85 2
262 248
262 248
1 0 4 0 0 0 0 22 0 0 86 2
251 239
251 239
1 0 26 0 0 0 0 21 0 0 87 2
238 230
238 230
1 0 27 0 0 0 0 20 0 0 88 2
220 221
220 221
1 0 28 0 0 0 0 19 0 0 89 2
201 212
201 212
1 0 29 0 0 0 0 18 0 0 90 2
179 203
179 203
1 0 30 0 0 0 0 17 0 0 91 2
158 194
158 194
8 0 3 0 0 128 0 43 0 0 0 2
270 257
258 257
7 0 3 0 0 128 0 43 0 0 0 2
270 248
250 248
6 0 4 0 0 128 0 43 0 0 0 2
270 239
236 239
5 0 26 0 0 4224 0 43 0 0 0 2
270 230
223 230
4 0 27 0 0 4224 0 43 0 0 0 2
270 221
205 221
3 0 28 0 0 4224 0 43 0 0 0 2
270 212
183 212
2 0 29 0 0 4224 0 43 0 0 0 2
270 203
161 203
1 0 30 0 0 4224 0 43 0 0 0 2
270 194
144 194
9 1 9 0 0 0 0 48 25 0 0 2
340 70
591 70
1 0 31 0 0 4096 0 46 0 0 101 2
545 152
545 133
1 0 32 0 0 0 0 47 0 0 102 2
545 124
545 124
1 0 6 0 0 0 0 26 0 0 98 2
469 97
469 97
1 0 7 0 0 0 0 27 0 0 99 2
492 88
492 88
1 0 8 0 0 0 0 28 0 0 100 2
516 79
516 79
12 0 6 0 0 0 0 48 0 0 0 2
334 97
489 97
11 0 7 0 0 0 0 48 0 0 0 2
334 88
511 88
10 0 8 0 0 0 0 48 0 0 0 2
334 79
532 79
14 0 31 0 0 4224 0 48 0 0 0 2
340 133
551 133
13 0 32 0 0 4224 0 48 0 0 0 2
334 124
550 124
1 0 4 0 0 0 0 29 0 0 111 2
267 133
267 133
1 0 4 0 0 0 0 30 0 0 112 2
262 124
262 124
1 0 33 0 0 0 0 31 0 0 113 2
251 115
251 115
1 0 34 0 0 0 0 32 0 0 114 2
238 106
238 106
1 0 35 0 0 0 0 33 0 0 115 2
220 97
220 97
1 0 36 0 0 0 0 34 0 0 116 2
201 88
201 88
1 0 37 0 0 0 0 35 0 0 117 2
179 79
179 79
1 0 38 0 0 0 0 36 0 0 118 2
158 70
158 70
8 0 4 0 0 128 0 48 0 0 0 2
270 133
258 133
7 0 4 0 0 128 0 48 0 0 0 2
270 124
250 124
6 0 33 0 0 4224 0 48 0 0 0 2
270 115
236 115
5 0 34 0 0 4224 0 48 0 0 0 2
270 106
223 106
4 0 35 0 0 4224 0 48 0 0 0 2
270 97
205 97
3 0 36 0 0 4224 0 48 0 0 0 2
270 88
183 88
2 0 37 0 0 4224 0 48 0 0 0 2
270 79
161 79
1 0 38 0 0 4224 0 48 0 0 0 2
270 70
144 70
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
