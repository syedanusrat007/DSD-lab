CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 129 583 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
3 V12
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
961 0 0
2
42920.9 0
0
13 Logic Switch~
5 174 568 0 1 11
0 19
0
0 0 21344 180
2 0V
-5 -16 9 -8
3 V11
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3178 0 0
2
42920.9 1
0
13 Logic Switch~
5 115 476 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
42920.9 2
0
13 Logic Switch~
5 103 151 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3951 0 0
2
42920.9 3
0
13 Logic Switch~
5 106 169 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
42920.9 4
0
13 Logic Switch~
5 381 66 0 1 11
0 15
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
42920.9 5
0
13 Logic Switch~
5 407 66 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 782
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9265 0 0
2
42920.9 6
0
13 Logic Switch~
5 431 66 0 1 11
0 13
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9442 0 0
2
42920.9 7
0
13 Logic Switch~
5 454 67 0 1 11
0 12
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
42920.9 8
0
13 Logic Switch~
5 114 503 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
42920.9 9
0
13 Logic Switch~
5 114 396 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9281 0 0
2
42920.9 10
0
13 Logic Switch~
5 113 289 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8464 0 0
2
42920.9 11
0
9 Inverter~
13 209 521 0 2 22
0 6 8
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
7168 0 0
2
42920.9 12
0
9 Inverter~
13 208 415 0 2 22
0 5 9
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3171 0 0
2
42920.9 13
0
9 Inverter~
13 190 307 0 2 22
0 4 10
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U5B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4139 0 0
2
42920.9 14
0
9 Inverter~
13 180 192 0 2 22
0 3 11
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6435 0 0
2
42920.9 15
0
7 74LS151
20 247 133 0 14 29
0 2 19 4 7 4 18 11 3 15
14 13 12 17 16
0
0 0 4832 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 1 0 0 0
1 U
5283 0 0
2
42920.9 16
0
14 Logic Display~
6 492 142 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
42920.9 17
0
14 Logic Display~
6 512 166 0 1 2
10 16
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
42920.9 18
0
14 Logic Display~
6 520 500 0 1 2
10 20
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
42920.9 19
0
14 Logic Display~
6 500 476 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
42920.9 20
0
7 74LS151
20 250 467 0 14 29
0 2 19 3 5 22 5 8 6 15
14 13 12 21 20
0
0 0 4832 0
7 74LS151
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 1 0 0 0
1 U
8402 0 0
2
42920.9 21
0
14 Logic Display~
6 520 393 0 1 2
10 23
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
42920.9 22
0
14 Logic Display~
6 500 369 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
42920.9 23
0
7 74LS151
20 250 360 0 14 29
0 2 19 6 4 6 4 9 5 15
14 13 12 24 23
0
0 0 4832 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 1 0 0 0
1 U
6118 0 0
2
42920.9 24
0
7 74LS151
20 249 253 0 14 29
0 2 19 5 3 5 3 10 4 15
14 13 12 26 25
0
0 0 4832 0
7 74LS151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
42920.9 25
0
14 Logic Display~
6 499 262 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
42920.9 26
0
14 Logic Display~
6 519 286 0 1 2
10 25
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
42920.9 27
0
82
0 0 2 0 0 4096 0 0 0 62 4 2
126 440
55 440
0 0 2 0 0 0 0 0 0 72 4 2
125 333
55 333
0 0 2 0 0 4096 0 0 0 82 4 2
130 226
55 226
0 1 2 0 0 8320 0 0 1 52 0 4
118 106
55 106
55 583
115 583
0 0 3 0 0 12416 0 0 0 45 60 6
143 169
143 91
14 91
14 548
145 548
145 458
0 0 4 0 0 4224 0 0 0 75 50 2
148 289
148 124
0 0 5 0 0 4224 0 0 0 65 80 2
154 396
154 244
0 0 6 0 0 4224 0 0 0 55 70 2
159 503
159 351
0 0 7 0 0 12416 0 0 0 0 49 6
173 506
173 525
38 525
38 82
208 82
208 133
0 0 5 0 0 0 0 0 0 65 59 2
166 396
166 467
0 0 4 0 0 0 0 0 0 75 69 2
169 289
169 360
0 0 3 0 0 0 0 0 0 45 79 2
198 169
198 253
0 0 4 0 0 0 0 0 0 75 48 2
159 289
159 142
0 0 5 0 0 0 0 0 0 65 78 2
176 396
176 262
0 0 6 0 0 0 0 0 0 55 68 2
182 503
182 369
0 0 5 0 0 0 0 0 0 65 57 2
187 396
187 485
0 0 4 0 0 0 0 0 0 75 67 2
209 289
209 378
0 0 3 0 0 0 0 0 0 45 77 2
209 169
209 271
2 0 8 0 0 8192 0 13 0 0 56 3
212 539
197 539
197 494
2 0 9 0 0 8192 0 14 0 0 66 3
211 433
196 433
196 387
2 0 10 0 0 8192 0 15 0 0 76 3
193 325
179 325
179 280
1 0 6 0 0 0 0 13 0 0 55 2
212 503
212 503
1 0 5 0 0 0 0 14 0 0 65 2
211 397
211 396
1 0 4 0 0 0 0 15 0 0 75 2
193 289
193 289
2 0 11 0 0 8192 0 16 0 0 46 3
183 210
167 210
167 160
1 0 3 0 0 0 0 16 0 0 45 2
183 174
183 169
12 0 12 0 0 8320 0 22 0 0 41 3
282 467
403 467
403 133
12 0 12 0 0 0 0 25 0 0 41 3
282 360
393 360
393 133
0 12 12 0 0 0 0 0 26 41 0 3
384 133
384 253
281 253
11 0 13 0 0 8320 0 22 0 0 42 3
282 458
375 458
375 124
0 11 13 0 0 0 0 0 25 42 0 3
364 124
364 351
282 351
11 0 13 0 0 0 0 26 0 0 42 3
281 244
356 244
356 124
0 10 14 0 0 4224 0 0 22 43 0 3
344 115
344 449
282 449
0 10 14 0 0 0 0 0 25 43 0 3
330 115
330 342
282 342
0 10 14 0 0 0 0 0 26 43 0 3
320 115
320 235
281 235
0 9 15 0 0 4224 0 0 22 44 0 3
310 106
310 440
288 440
0 9 15 0 0 0 0 0 25 44 0 3
301 106
301 333
288 333
0 9 15 0 0 0 0 0 26 44 0 3
290 106
290 226
287 226
14 1 16 0 0 4224 0 17 19 0 0 2
285 169
497 169
13 1 17 0 0 4224 0 17 18 0 0 2
279 160
492 160
12 1 12 0 0 0 0 17 9 0 0 4
279 133
455 133
455 79
454 79
11 1 13 0 0 0 0 17 8 0 0 3
279 124
431 124
431 78
10 1 14 0 0 0 0 17 7 0 0 3
279 115
407 115
407 78
9 1 15 0 0 0 0 17 6 0 0 3
285 106
381 106
381 78
8 1 3 0 0 0 0 17 5 0 0 2
215 169
118 169
7 0 11 0 0 4224 0 17 0 0 0 2
215 160
114 160
6 1 18 0 0 4224 0 17 4 0 0 2
215 151
115 151
5 0 4 0 0 0 0 17 0 0 0 2
215 142
118 142
4 0 7 0 0 0 0 17 0 0 0 2
215 133
116 133
3 0 4 0 0 0 0 17 0 0 0 2
215 124
114 124
2 1 19 0 0 8320 0 17 2 0 0 4
215 115
78 115
78 568
160 568
1 0 2 0 0 0 0 17 0 0 0 2
215 106
114 106
14 1 20 0 0 4224 0 22 20 0 0 2
288 503
505 503
13 1 21 0 0 4224 0 22 21 0 0 2
282 494
500 494
8 1 6 0 0 0 0 22 10 0 0 2
218 503
126 503
7 0 8 0 0 4224 0 22 0 0 0 2
218 494
122 494
6 0 5 0 0 0 0 22 0 0 0 2
218 485
123 485
5 1 22 0 0 4224 0 22 3 0 0 2
218 476
127 476
4 0 5 0 0 0 0 22 0 0 0 2
218 467
124 467
3 0 3 0 0 0 0 22 0 0 0 2
218 458
122 458
2 0 19 0 0 0 0 22 0 0 51 2
218 449
78 449
1 0 2 0 0 0 0 22 0 0 0 2
218 440
122 440
14 1 23 0 0 4224 0 25 23 0 0 2
288 396
505 396
13 1 24 0 0 4224 0 25 24 0 0 2
282 387
500 387
8 1 5 0 0 0 0 25 11 0 0 2
218 396
126 396
7 0 9 0 0 4224 0 25 0 0 0 2
218 387
122 387
6 0 4 0 0 0 0 25 0 0 0 2
218 378
123 378
5 0 6 0 0 0 0 25 0 0 0 2
218 369
126 369
4 0 4 0 0 0 0 25 0 0 0 2
218 360
124 360
3 0 6 0 0 0 0 25 0 0 0 2
218 351
122 351
2 0 19 0 0 0 0 25 0 0 51 2
218 342
78 342
1 0 2 0 0 0 0 25 0 0 0 2
218 333
122 333
14 1 25 0 0 4224 0 26 28 0 0 2
287 289
504 289
13 1 26 0 0 4224 0 26 27 0 0 2
281 280
499 280
8 1 4 0 0 0 0 26 12 0 0 2
217 289
125 289
7 0 10 0 0 4224 0 26 0 0 0 2
217 280
121 280
6 0 3 0 0 0 0 26 0 0 0 2
217 271
122 271
5 0 5 0 0 0 0 26 0 0 0 2
217 262
125 262
4 0 3 0 0 0 0 26 0 0 0 2
217 253
123 253
3 0 5 0 0 0 0 26 0 0 0 2
217 244
121 244
2 0 19 0 0 0 0 26 0 0 51 2
217 235
78 235
1 0 2 0 0 0 0 26 0 0 0 2
217 226
121 226
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
