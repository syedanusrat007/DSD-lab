CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
75
13 Logic Switch~
5 866 1044 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
3 V13
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7788 0 0
2
5.89808e-315 0
0
13 Logic Switch~
5 661 55 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
3 V12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3273 0 0
2
5.89808e-315 0
0
13 Logic Switch~
5 598 54 0 1 11
0 54
0
0 0 21360 782
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3761 0 0
2
5.89808e-315 5.26354e-315
0
13 Logic Switch~
5 533 53 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3226 0 0
2
5.89808e-315 5.30499e-315
0
13 Logic Switch~
5 480 52 0 1 11
0 25
0
0 0 21360 782
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4244 0 0
2
5.89808e-315 5.32571e-315
0
13 Logic Switch~
5 427 56 0 1 11
0 66
0
0 0 21360 782
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5225 0 0
2
5.89808e-315 5.34643e-315
0
13 Logic Switch~
5 370 54 0 10 11
0 55 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
768 0 0
2
5.89808e-315 5.3568e-315
0
13 Logic Switch~
5 317 52 0 1 11
0 41
0
0 0 21360 782
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5735 0 0
2
5.89808e-315 5.36716e-315
0
13 Logic Switch~
5 271 54 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5881 0 0
2
5.89808e-315 5.37752e-315
0
13 Logic Switch~
5 202 53 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3275 0 0
2
5.89808e-315 5.38788e-315
0
13 Logic Switch~
5 139 53 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4203 0 0
2
5.89808e-315 5.39306e-315
0
13 Logic Switch~
5 73 52 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
5.89808e-315 5.39824e-315
0
13 Logic Switch~
5 19 57 0 1 11
0 9
0
0 0 21360 782
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9102 0 0
2
5.89808e-315 5.40342e-315
0
9 2-In XOR~
219 893 1035 0 3 22
0 3 2 60
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U16D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
5586 0 0
2
5.89808e-315 0
0
9 2-In XOR~
219 845 1026 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U16C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
525 0 0
2
5.89808e-315 0
0
9 4-In NOR~
219 778 1055 0 5 22
0 68 69 6 7 4
0
0 0 624 692
4 4002
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 1 19 0
1 U
6206 0 0
2
5.89808e-315 0
0
9 2-In XOR~
219 755 1014 0 3 22
0 7 6 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U16B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
3418 0 0
2
5.89808e-315 0
0
9 2-In AND~
219 916 1138 0 3 22
0 11 9 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
9312 0 0
2
5.89808e-315 0
0
9 4-In NOR~
219 822 1129 0 5 22
0 70 71 8 12 11
0
0 0 624 692
4 4002
-14 -24 14 -16
4 U17B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 2 18 0
1 U
7419 0 0
2
5.89808e-315 0
0
14 Logic Display~
6 2024 115 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
472 0 0
2
5.89808e-315 5.4086e-315
0
14 Logic Display~
6 1961 123 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4714 0 0
2
5.89808e-315 5.41378e-315
0
14 Logic Display~
6 1877 114 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9386 0 0
2
5.89808e-315 5.41896e-315
0
9 4-In NOR~
219 1871 164 0 5 22
0 14 17 16 15 18
0
0 0 624 90
4 4002
-14 -24 14 -16
4 U17A
30 -2 58 6
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 18 0
1 U
7610 0 0
2
5.89808e-315 5.42414e-315
0
14 Logic Display~
6 1768 122 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
5.89808e-315 5.42933e-315
0
9 2-In XOR~
219 1765 167 0 3 22
0 19 13 20
0
0 0 624 602
6 74LS86
-21 -24 21 -16
4 U16A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
3608 0 0
2
5.89808e-315 5.43192e-315
0
14 Logic Display~
6 1647 106 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6397 0 0
2
5.89808e-315 5.43451e-315
0
14 Logic Display~
6 1608 107 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3967 0 0
2
5.89808e-315 5.4371e-315
0
14 Logic Display~
6 1573 107 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8621 0 0
2
5.89808e-315 5.43969e-315
0
14 Logic Display~
6 1446 111 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89808e-315 5.44228e-315
0
14 Logic Display~
6 1526 109 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7385 0 0
2
5.89808e-315 5.44487e-315
0
8 2-In OR~
219 1322 961 0 3 22
0 50 49 40
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
6519 0 0
2
5.89808e-315 5.44746e-315
0
9 Inverter~
13 675 70 0 2 22
0 65 64
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 15 0
1 U
552 0 0
2
5.89808e-315 5.45005e-315
0
9 Inverter~
13 611 71 0 2 22
0 54 53
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 15 0
1 U
5551 0 0
2
5.89808e-315 5.45264e-315
0
9 Inverter~
13 547 70 0 2 22
0 45 44
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 15 0
1 U
8715 0 0
2
5.89808e-315 5.45523e-315
0
9 Inverter~
13 495 69 0 2 22
0 25 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 15 0
1 U
9763 0 0
2
5.89808e-315 5.45782e-315
0
9 Inverter~
13 153 69 0 2 22
0 8 67
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 15 0
1 U
8443 0 0
2
5.89808e-315 5.46041e-315
0
9 Inverter~
13 32 72 0 2 22
0 9 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 15 0
1 U
3719 0 0
2
5.89808e-315 5.463e-315
0
8 2-In OR~
219 1013 190 0 3 22
0 10 33 31
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8671 0 0
2
5.89808e-315 5.47077e-315
0
9 2-In AND~
219 904 305 0 3 22
0 8 25 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7168 0 0
2
5.89808e-315 5.47207e-315
0
9 2-In AND~
219 905 346 0 3 22
0 12 24 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
49 0 0
2
5.89808e-315 5.47336e-315
0
8 2-In OR~
219 959 322 0 3 22
0 27 26 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6536 0 0
2
5.89808e-315 5.47466e-315
0
9 2-In XOR~
219 1189 211 0 3 22
0 31 30 32
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3931 0 0
2
5.89808e-315 5.47595e-315
0
9 2-In XOR~
219 1187 274 0 3 22
0 22 32 14
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4390 0 0
2
5.89808e-315 5.47725e-315
0
9 2-In AND~
219 1191 141 0 3 22
0 19 7 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3242 0 0
2
5.89808e-315 5.47854e-315
0
9 2-In AND~
219 1260 311 0 3 22
0 22 32 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6760 0 0
2
5.89808e-315 5.47984e-315
0
9 2-In AND~
219 1264 358 0 3 22
0 31 30 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5760 0 0
2
5.89808e-315 5.48113e-315
0
8 2-In OR~
219 1320 331 0 3 22
0 29 28 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3781 0 0
2
5.89808e-315 5.48243e-315
0
8 2-In OR~
219 1324 636 0 3 22
0 34 35 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8545 0 0
2
5.89808e-315 5.48372e-315
0
9 2-In AND~
219 1268 663 0 3 22
0 37 36 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9739 0 0
2
5.89808e-315 5.48502e-315
0
9 2-In AND~
219 1264 616 0 3 22
0 39 38 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
388 0 0
2
5.89808e-315 5.48631e-315
0
9 2-In AND~
219 1195 446 0 3 22
0 40 7 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
4595 0 0
2
5.89808e-315 5.48761e-315
0
9 2-In XOR~
219 1191 579 0 3 22
0 39 38 17
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3173 0 0
2
5.89808e-315 5.4889e-315
0
9 2-In XOR~
219 1193 516 0 3 22
0 37 36 39
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9261 0 0
2
5.89808e-315 5.4902e-315
0
8 2-In OR~
219 963 627 0 3 22
0 43 42 36
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-4 -28 17 -20
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3494 0 0
2
5.89808e-315 5.49149e-315
0
9 2-In AND~
219 909 651 0 3 22
0 12 44 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9101 0 0
2
5.89808e-315 5.49279e-315
0
9 2-In AND~
219 908 610 0 3 22
0 8 45 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
358 0 0
2
5.89808e-315 5.49408e-315
0
8 2-In OR~
219 1019 493 0 3 22
0 10 41 37
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3726 0 0
2
5.89808e-315 5.49538e-315
0
9 2-In AND~
219 1267 988 0 3 22
0 47 46 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
999 0 0
2
5.89808e-315 5.49926e-315
0
9 2-In AND~
219 1263 941 0 3 22
0 48 23 50
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
8787 0 0
2
5.89808e-315 5.50056e-315
0
9 2-In AND~
219 1184 760 0 3 22
0 56 7 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3348 0 0
2
5.89808e-315 5.50185e-315
0
9 2-In XOR~
219 1190 904 0 3 22
0 48 23 16
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3395 0 0
2
5.89808e-315 5.50315e-315
0
9 2-In XOR~
219 1192 841 0 3 22
0 47 46 48
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
7740 0 0
2
5.89808e-315 5.50444e-315
0
8 2-In OR~
219 962 952 0 3 22
0 52 51 46
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
6480 0 0
2
5.89808e-315 5.50574e-315
0
9 2-In AND~
219 908 976 0 3 22
0 12 53 51
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
342 0 0
2
5.89808e-315 5.50703e-315
0
9 2-In AND~
219 907 935 0 3 22
0 8 54 52
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
9953 0 0
2
5.89808e-315 5.50833e-315
0
8 2-In OR~
219 1016 820 0 3 22
0 10 55 47
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
361 0 0
2
5.89808e-315 5.50963e-315
0
8 2-In OR~
219 1328 1291 0 3 22
0 58 57 56
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3343 0 0
2
5.89808e-315 5.51286e-315
0
9 2-In AND~
219 1272 1318 0 3 22
0 21 59 57
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
7923 0 0
2
5.89808e-315 5.51351e-315
0
9 2-In AND~
219 1279 1273 0 3 22
0 61 60 58
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
6174 0 0
2
5.89808e-315 5.51416e-315
0
9 2-In XOR~
219 1195 1234 0 3 22
0 61 60 15
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
6692 0 0
2
5.89808e-315 5.51545e-315
0
9 2-In XOR~
219 1197 1171 0 3 22
0 21 59 61
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
8790 0 0
2
5.89808e-315 5.5161e-315
0
8 2-In OR~
219 967 1282 0 3 22
0 63 62 59
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4595 0 0
2
5.89808e-315 5.51675e-315
0
9 2-In AND~
219 913 1306 0 3 22
0 12 64 62
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
667 0 0
2
5.89808e-315 5.5174e-315
0
9 2-In AND~
219 912 1265 0 3 22
0 8 65 63
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
8743 0 0
2
5.89808e-315 5.51804e-315
0
8 2-In OR~
219 1021 1150 0 3 22
0 10 66 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
8298 0 0
2
5.89808e-315 5.51869e-315
0
134
1 2 2 0 0 4224 0 1 14 0 0 2
878 1044
877 1044
1 3 3 0 0 4224 0 14 15 0 0 2
877 1026
878 1026
5 2 4 0 0 4224 0 16 15 0 0 3
817 1055
817 1035
829 1035
3 1 5 0 0 8320 0 17 15 0 0 3
788 1014
788 1017
829 1017
0 3 6 0 0 8192 0 0 16 7 0 3
708 1023
708 1050
761 1050
0 4 7 0 0 8192 0 0 16 8 0 3
722 1005
722 1041
761 1041
2 0 6 0 0 4096 0 17 0 0 131 2
739 1023
202 1023
1 0 7 0 0 4096 0 17 0 0 116 2
739 1005
53 1005
3 0 8 0 0 4096 0 19 0 0 132 2
805 1124
139 1124
2 0 9 0 0 8192 0 18 0 0 15 3
892 1147
892 1148
879 1148
1 0 10 0 0 4096 0 66 0 0 13 2
1003 811
994 811
1 0 10 0 0 4096 0 57 0 0 13 2
1006 484
994 484
0 1 10 0 0 4224 0 0 38 14 0 3
994 1141
994 181
1000 181
3 1 10 0 0 0 0 18 75 0 0 4
937 1138
936 1138
936 1141
1008 1141
0 0 9 0 0 12288 0 0 0 0 134 4
887 1148
829 1148
829 1174
19 1174
1 5 11 0 0 4224 0 18 19 0 0 2
892 1129
861 1129
4 0 12 0 0 12288 0 19 0 0 133 4
805 1115
789 1115
789 1106
73 1106
0 1 13 0 0 4224 0 0 20 41 0 3
1446 318
2024 318
2024 133
0 1 14 0 0 4096 0 0 21 23 0 3
1864 204
1961 204
1961 141
0 4 15 0 0 4096 0 0 23 32 0 3
1647 302
1891 302
1891 187
0 3 16 0 0 4096 0 0 23 33 0 3
1608 283
1882 283
1882 187
0 2 17 0 0 4096 0 0 23 34 0 3
1573 259
1873 259
1873 187
0 1 14 0 0 4224 0 0 23 47 0 3
1526 239
1864 239
1864 187
1 5 18 0 0 4224 0 22 23 0 0 2
1877 132
1877 131
0 1 19 0 0 4096 0 0 25 54 0 3
1390 217
1777 217
1777 186
2 0 13 0 0 0 0 25 0 0 41 2
1759 186
1446 186
1 3 20 0 0 4224 0 24 25 0 0 2
1768 140
1768 137
1 0 21 0 0 8320 0 68 0 0 29 3
1248 1309
1153 1309
1153 1162
1 3 21 0 0 0 0 71 75 0 0 4
1181 1162
1070 1162
1070 1150
1054 1150
0 1 22 0 0 8192 0 0 45 49 0 3
1160 265
1160 302
1236 302
0 2 23 0 0 8192 0 0 59 81 0 3
1167 913
1167 950
1239 950
1 3 15 0 0 4224 0 26 70 0 0 3
1647 124
1647 1234
1228 1234
1 3 16 0 0 4224 0 27 61 0 0 3
1608 125
1608 904
1223 904
1 3 17 0 0 4224 0 28 52 0 0 3
1573 125
1573 579
1224 579
2 0 24 0 0 4096 0 40 0 0 114 2
881 355
516 355
1 0 12 0 0 4096 0 40 0 0 133 2
881 337
73 337
2 0 25 0 0 4096 0 39 0 0 126 2
880 314
480 314
1 0 8 0 0 4096 0 39 0 0 132 2
880 296
139 296
3 2 26 0 0 8320 0 40 41 0 0 4
926 346
933 346
933 331
946 331
3 1 27 0 0 4224 0 39 41 0 0 4
925 305
937 305
937 313
946 313
3 1 13 0 0 0 0 47 29 0 0 3
1353 331
1446 331
1446 129
3 2 28 0 0 8320 0 46 47 0 0 4
1285 358
1296 358
1296 340
1307 340
3 1 29 0 0 8320 0 45 47 0 0 3
1281 311
1281 322
1307 322
2 0 30 0 0 4224 0 46 0 0 50 3
1240 367
1048 367
1048 322
1 0 31 0 0 8320 0 46 0 0 51 3
1240 349
1103 349
1103 190
0 2 32 0 0 8192 0 0 45 48 0 3
1154 283
1154 320
1236 320
3 1 14 0 0 0 0 43 30 0 0 3
1220 274
1526 274
1526 127
3 2 32 0 0 12416 0 42 43 0 0 6
1222 211
1323 211
1323 241
1112 241
1112 283
1171 283
3 1 22 0 0 12416 0 44 43 0 0 6
1212 141
1323 141
1323 176
1131 176
1131 265
1171 265
3 2 30 0 0 0 0 41 42 0 0 4
992 322
1081 322
1081 220
1173 220
3 1 31 0 0 0 0 38 42 0 0 4
1046 190
1152 190
1152 202
1173 202
2 0 7 0 0 4096 0 44 0 0 116 2
1167 150
53 150
2 0 33 0 0 12288 0 38 0 0 130 4
1000 199
938 199
938 234
271 234
0 1 19 0 0 4224 0 0 44 55 0 5
1390 636
1390 94
1119 94
1119 132
1167 132
3 0 19 0 0 0 0 48 0 0 0 2
1357 636
1515 636
3 1 34 0 0 8320 0 50 48 0 0 3
1285 616
1285 627
1311 627
3 2 35 0 0 8320 0 49 48 0 0 4
1289 663
1298 663
1298 645
1311 645
2 0 36 0 0 4224 0 49 0 0 66 3
1244 672
1066 672
1066 627
1 0 37 0 0 8320 0 49 0 0 67 3
1244 654
1099 654
1099 493
0 2 38 0 0 8192 0 0 50 64 0 3
1171 588
1171 625
1240 625
0 1 39 0 0 4096 0 0 50 65 0 3
1233 516
1233 607
1240 607
2 0 7 0 0 4096 0 51 0 0 116 2
1171 455
53 455
0 1 40 0 0 4224 0 0 51 80 0 5
1370 961
1370 409
1147 409
1147 437
1171 437
3 2 38 0 0 12416 0 51 52 0 0 6
1216 446
1259 446
1259 478
1115 478
1115 588
1175 588
3 1 39 0 0 12416 0 53 52 0 0 6
1226 516
1293 516
1293 542
1125 542
1125 570
1175 570
3 2 36 0 0 0 0 54 53 0 0 4
996 627
1076 627
1076 525
1177 525
3 1 37 0 0 0 0 57 53 0 0 4
1052 493
1143 493
1143 507
1177 507
0 2 41 0 0 4096 0 0 57 129 0 4
317 530
985 530
985 502
1006 502
3 2 42 0 0 8320 0 55 54 0 0 3
930 651
930 636
950 636
3 1 43 0 0 8320 0 56 54 0 0 3
929 610
929 618
950 618
2 0 44 0 0 4096 0 55 0 0 113 2
885 660
568 660
1 0 12 0 0 4096 0 55 0 0 133 2
885 642
73 642
2 0 45 0 0 4096 0 56 0 0 125 2
884 619
533 619
1 0 8 0 0 4096 0 56 0 0 132 2
884 601
139 601
2 0 46 0 0 4224 0 58 0 0 83 3
1243 997
1099 997
1099 952
1 0 47 0 0 8320 0 58 0 0 84 3
1243 979
1158 979
1158 832
0 1 48 0 0 4096 0 0 59 82 0 3
1230 841
1230 932
1239 932
3 2 49 0 0 8320 0 58 31 0 0 3
1288 988
1288 970
1309 970
3 1 50 0 0 8320 0 59 31 0 0 3
1284 941
1284 952
1309 952
3 0 40 0 0 0 0 31 0 0 0 2
1355 961
1510 961
3 2 23 0 0 12416 0 60 61 0 0 6
1205 760
1266 760
1266 810
1089 810
1089 913
1174 913
3 1 48 0 0 12416 0 62 61 0 0 6
1225 841
1281 841
1281 869
1160 869
1160 895
1174 895
3 2 46 0 0 0 0 63 62 0 0 4
995 952
1125 952
1125 850
1176 850
3 1 47 0 0 0 0 66 62 0 0 4
1049 820
1132 820
1132 832
1176 832
2 0 7 0 0 0 0 60 0 0 116 2
1160 769
53 769
3 2 51 0 0 8320 0 64 63 0 0 4
929 976
936 976
936 961
949 961
3 1 52 0 0 8320 0 65 63 0 0 4
928 935
928 946
949 946
949 943
2 0 53 0 0 4096 0 64 0 0 112 2
884 985
632 985
1 0 12 0 0 0 0 64 0 0 133 2
884 967
73 967
2 0 54 0 0 4096 0 65 0 0 124 2
883 944
598 944
1 0 8 0 0 0 0 65 0 0 132 2
883 926
139 926
2 0 55 0 0 12288 0 66 0 0 128 4
1003 829
983 829
983 862
370 862
0 1 56 0 0 4224 0 0 60 94 0 5
1399 1291
1399 731
1157 731
1157 751
1160 751
3 0 56 0 0 0 0 67 0 0 0 2
1361 1291
1557 1291
3 2 57 0 0 8320 0 68 67 0 0 4
1293 1318
1304 1318
1304 1300
1315 1300
3 1 58 0 0 8320 0 69 67 0 0 3
1300 1273
1300 1282
1315 1282
2 0 59 0 0 8320 0 68 0 0 103 3
1248 1327
1170 1327
1170 1180
2 0 60 0 0 4096 0 69 0 0 100 3
1255 1282
1115 1282
1115 1243
0 1 61 0 0 4096 0 0 69 102 0 5
1256 1171
1256 1243
1230 1243
1230 1264
1255 1264
3 2 60 0 0 16512 0 14 70 0 0 6
926 1035
927 1035
927 1040
1106 1040
1106 1243
1179 1243
1 0 61 0 0 12416 0 70 0 0 102 5
1179 1225
1132 1225
1132 1201
1240 1201
1240 1171
3 0 61 0 0 0 0 71 0 0 0 2
1230 1171
1279 1171
3 2 59 0 0 0 0 72 71 0 0 4
1000 1282
1076 1282
1076 1180
1181 1180
3 2 62 0 0 8320 0 73 72 0 0 3
934 1306
934 1291
954 1291
3 1 63 0 0 8320 0 74 72 0 0 3
933 1265
933 1273
954 1273
1 0 12 0 0 4096 0 73 0 0 133 2
889 1297
73 1297
2 0 64 0 0 4096 0 73 0 0 111 2
889 1315
696 1315
2 0 65 0 0 4096 0 74 0 0 123 2
888 1274
661 1274
1 0 8 0 0 4096 0 74 0 0 132 2
888 1256
139 1256
2 0 66 0 0 12288 0 75 0 0 127 4
1008 1159
953 1159
953 1188
427 1188
2 0 64 0 0 4224 0 32 0 0 0 2
696 70
696 1373
2 0 53 0 0 4224 0 33 0 0 0 2
632 71
632 1373
2 0 44 0 0 4224 0 34 0 0 0 2
568 70
568 1372
2 0 24 0 0 4224 0 35 0 0 0 2
516 69
516 1371
2 0 67 0 0 4224 0 36 0 0 0 2
174 69
174 1364
2 0 7 0 0 4224 0 37 0 0 0 2
53 72
53 1358
1 0 65 0 0 0 0 32 0 0 123 2
660 70
661 70
1 0 54 0 0 0 0 33 0 0 124 2
596 71
598 71
1 0 45 0 0 0 0 34 0 0 125 2
532 70
533 70
1 0 25 0 0 0 0 35 0 0 126 2
480 69
480 69
1 0 8 0 0 0 0 36 0 0 132 2
138 69
139 69
1 0 9 0 0 0 0 37 0 0 134 2
17 72
19 72
1 0 65 0 0 4224 0 2 0 0 0 2
661 67
661 1367
1 0 54 0 0 4224 0 3 0 0 0 2
598 66
598 1369
1 0 45 0 0 4224 0 4 0 0 0 2
533 65
533 1370
1 0 25 0 0 4224 0 5 0 0 0 2
480 64
480 1369
1 0 66 0 0 4224 0 6 0 0 0 2
427 68
427 1369
1 0 55 0 0 4224 0 7 0 0 0 2
370 66
370 1371
1 0 41 0 0 4224 0 8 0 0 0 2
317 64
317 1373
1 0 33 0 0 4224 0 9 0 0 0 2
271 66
271 1370
1 0 6 0 0 4224 0 10 0 0 0 2
202 65
202 1368
1 0 8 0 0 4224 0 11 0 0 0 2
139 65
139 1364
1 0 12 0 0 4224 0 12 0 0 0 2
73 64
73 1359
1 0 9 0 0 4224 0 13 0 0 0 2
19 69
19 1361
68
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 17
840 1161 1010 1192
847 1165 1002 1186
17 (s1 nor s0)and s2
-16 0 0 0 400 255 0 0 0 3 2 1 18
12 Cooper Black
0 0 0 9
800 1083 891 1110
808 1087 882 1106
9 s1 nor s0
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
950 1009 990 1036
957 1013 982 1032
2 z1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1210 728 1250 755
1217 732 1242 751
2 z2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1210 410 1250 437
1217 414 1242 433
2 z3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1205 100 1245 127
1212 104 1237 123
2 z4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1349 299 1384 326
1353 303 1379 322
2 c5
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1349 605 1384 632
1353 609 1379 628
2 c4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1356 930 1391 957
1360 934 1386 953
2 c3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1357 1261 1398 1288
1364 1265 1390 1284
2 c2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
998 1253 1041 1280
1005 1257 1033 1276
2 y1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1051 1121 1094 1148
1058 1125 1086 1144
2 x1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
984 912 1027 939
991 916 1019 935
2 y2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1037 780 1080 807
1044 784 1072 803
2 x2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
993 599 1036 626
1000 603 1028 622
2 y3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1043 464 1086 491
1050 468 1078 487
2 x3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
983 282 1024 309
989 286 1017 305
2 y4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1217 240 1251 267
1221 244 1246 263
2 f4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1225 547 1259 574
1229 551 1254 570
2 f3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1223 874 1257 901
1227 878 1252 897
2 f2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1226 1201 1260 1228
1230 1205 1255 1224
2 f1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1037 152 1074 179
1041 156 1069 175
2 x4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1 1 40 28
8 5 32 24
2 s2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
58 0 97 27
65 4 89 23
2 s1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
125 1 164 28
132 5 156 24
2 s0
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
188 2 229 29
195 6 221 25
2 c1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
254 3 295 30
261 7 287 26
2 a4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
303 1 344 28
310 5 336 24
2 a3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
358 3 399 30
365 7 391 26
2 a2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
412 4 453 31
419 8 445 27
2 a1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
463 2 504 29
470 6 496 25
2 b4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
517 3 558 30
524 7 550 26
2 b3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
580 3 621 30
587 7 613 26
2 b2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
643 4 684 31
650 8 676 27
2 b1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
658 1371 699 1398
665 1375 691 1394
2 b1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
595 1372 636 1399
602 1376 628 1395
2 b2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
530 1372 571 1399
537 1376 563 1395
2 b3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
480 1370 521 1397
487 1374 513 1393
2 b4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
419 1376 460 1403
426 1380 452 1399
2 a1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
365 1375 406 1402
372 1379 398 1398
2 a2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
310 1373 351 1400
317 1377 343 1396
2 a3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
183 1368 224 1395
190 1372 216 1391
2 c1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
136 1367 175 1394
143 1371 167 1390
2 s0
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
54 1358 93 1385
61 1362 85 1381
2 s1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
12 1362 51 1389
19 1366 43 1385
2 s2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
258 1371 293 1398
262 1375 288 1394
2 a4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
659 546 700 573
666 550 692 569
2 b1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
595 546 636 573
602 550 628 569
2 b2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
531 545 572 572
538 549 564 568
2 b3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
477 546 518 573
484 550 510 569
2 b4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
431 548 472 575
438 552 464 571
2 a1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
370 543 411 570
377 547 403 566
2 a2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
313 543 354 570
320 547 346 566
2 a3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
269 542 310 569
276 546 302 565
2 a4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
198 544 239 571
205 548 231 567
2 c1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
136 548 175 575
143 552 167 571
2 s0
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
69 547 108 574
76 551 100 570
2 s1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
15 547 54 574
22 551 46 570
2 s2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1425 56 1466 83
1432 60 1458 79
2 c5
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1505 54 1545 81
1512 58 1537 77
2 f4
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1548 53 1588 80
1555 57 1580 76
2 f3
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1586 55 1626 82
1593 59 1618 78
2 f2
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 2
1628 56 1668 83
1635 60 1660 79
2 f1
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 1
1752 63 1782 90
1759 67 1774 86
1 v
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 1
1862 62 1891 89
1869 66 1883 85
1 z
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 1
1945 62 1973 89
1952 66 1965 85
1 s
-16 0 0 0 700 0 0 0 0 3 2 1 18
12 Engravers MT
0 0 0 1
2009 55 2039 82
2016 59 2031 78
1 c
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 38
904 1042 1074 1099
911 1046 1066 1088
38 (((s2' xor c1)xor
(s2'nor c1)))xor 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
