CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 1970 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
181
13 Logic Switch~
5 1714 227 0 10 11
0 61 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3494 0 0
2
5.89774e-315 0
0
13 Logic Switch~
5 1147 217 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3507 0 0
2
42661 0
0
13 Logic Switch~
5 1786 296 0 10 11
0 89 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 CLR
-20 -18 1 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5151 0 0
2
42661 1
0
13 Logic Switch~
5 205 2033 0 1 11
0 100
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 SU
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3701 0 0
2
42661 2
0
13 Logic Switch~
5 202 2293 0 10 11
0 109 0 0 0 0 0 0 0 0
1
0
0 0 21232 0
2 5V
-6 -16 8 -8
2 C0
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8585 0 0
2
42661 3
0
13 Logic Switch~
5 204 2247 0 10 11
0 110 0 0 0 0 0 0 0 0
1
0
0 0 29424 0
2 5V
-6 -16 8 -8
2 C1
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8809 0 0
2
42661 4
0
13 Logic Switch~
5 204 2203 0 1 11
0 111
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 C2
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5993 0 0
2
42661 5
0
13 Logic Switch~
5 204 2158 0 1 11
0 112
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 C3
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8654 0 0
2
42661 6
0
13 Logic Switch~
5 211 1888 0 10 11
0 113 0 0 0 0 0 0 0 0
1
0
0 0 21232 0
2 5V
-6 -16 8 -8
2 B0
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7223 0 0
2
42661 7
0
13 Logic Switch~
5 210 1850 0 1 11
0 114
0
0 0 21232 0
2 0V
-6 -16 8 -8
2 B1
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3641 0 0
2
42661 8
0
13 Logic Switch~
5 211 1813 0 1 11
0 115
0
0 0 21232 0
2 0V
-6 -16 8 -8
2 B2
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3104 0 0
2
42661 9
0
13 Logic Switch~
5 210 1772 0 1 11
0 116
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 B3
-5 -22 9 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3296 0 0
2
42661 10
0
13 Logic Switch~
5 198 1416 0 10 11
0 117 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
3 EA6
-8 -22 13 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8534 0 0
2
42661 11
0
13 Logic Switch~
5 196 1389 0 1 11
0 118
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 EA5
-8 -22 13 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
949 0 0
2
42661 12
0
13 Logic Switch~
5 256 1489 0 10 11
0 119 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
3 EA4
-8 -22 13 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3371 0 0
2
42661 13
0
13 Logic Switch~
5 256 1464 0 1 11
0 120
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 EA3
-8 -22 13 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7311 0 0
2
42661 14
0
13 Logic Switch~
5 258 1439 0 1 11
0 121
0
0 0 20720 0
2 0V
-6 -16 8 -8
3 EA2
-8 -22 13 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
42661 15
0
13 Logic Switch~
5 258 1414 0 10 11
0 122 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
3 EA1
-8 -22 13 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3526 0 0
2
42661 16
0
13 Logic Switch~
5 267 710 0 1 11
0 133
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4129 0 0
2
42661 17
0
13 Logic Switch~
5 270 656 0 1 11
0 134
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6278 0 0
2
42661 18
0
13 Logic Switch~
5 270 607 0 1 11
0 135
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 A1
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3482 0 0
2
42661 19
0
13 Logic Switch~
5 272 557 0 1 11
0 136
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8323 0 0
2
42661 20
0
13 Logic Switch~
5 215 536 0 1 11
0 137
0
0 0 21360 0
2 0V
-6 -16 8 -8
7 SELECT1
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3984 0 0
2
42661 21
0
13 Logic Switch~
5 93 71 0 10 11
0 143 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7622 0 0
2
42661 22
0
8 3-In OR~
219 2550 822 0 4 22
0 7 6 5 4
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U14C
-2 23 26 31
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 10 0
1 U
816 0 0
2
42661.1 0
0
5 4071~
219 2376 1020 0 3 22
0 9 10 8
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U18C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 14 0
1 U
4656 0 0
2
42661.1 0
0
5 4081~
219 2253 828 0 3 22
0 13 12 11
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 15 0
1 U
6356 0 0
2
42661.1 0
0
5 4071~
219 2207 1003 0 3 22
0 15 16 14
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U18B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
7479 0 0
2
42661.1 0
0
8 4-In OR~
219 2179 931 0 5 22
0 7 6 5 17 15
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U16B
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 11 0
1 U
5690 0 0
2
42661.1 0
0
5 4081~
219 2142 851 0 3 22
0 13 18 17
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 15 0
1 U
5617 0 0
2
42661.1 0
0
5 4081~
219 2140 793 0 3 22
0 13 19 5
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19B
-31 -25 -3 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 15 0
1 U
3903 0 0
2
42661.1 0
0
5 4081~
219 2151 746 0 3 22
0 13 20 6
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
4452 0 0
2
42661.1 0
0
5 4081~
219 2141 679 0 3 22
0 13 21 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 13 0
1 U
6282 0 0
2
42661.1 0
0
8 3-In OR~
219 2094 1011 0 4 22
0 23 9 10 22
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U14B
-2 23 26 31
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
7187 0 0
2
42661.1 0
0
5 4081~
219 2055 976 0 3 22
0 13 24 10
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 13 0
1 U
6866 0 0
2
42661.1 0
0
5 4081~
219 2078 909 0 3 22
0 13 25 9
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U17B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 13 0
1 U
7670 0 0
2
42661.1 0
0
5 4071~
219 1954 722 0 3 22
0 16 28 29
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U18A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
951 0 0
2
42661.1 0
0
5 4081~
219 1948 649 0 3 22
0 32 31 16
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U17A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
9536 0 0
2
42661.1 0
0
8 4-In OR~
219 1883 619 0 5 22
0 30 23 34 26 33
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 11 0
1 U
5495 0 0
2
42661.1 0
0
5 4081~
219 1830 602 0 3 22
0 13 31 23
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 9 0
1 U
8152 0 0
2
42661.1 0
0
8 3-In OR~
219 1776 667 0 4 22
0 34 30 26 27
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U14A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
6223 0 0
2
42661.1 0
0
5 4081~
219 1693 696 0 3 22
0 32 25 26
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
5441 0 0
2
42661.1 0
0
5 4081~
219 1686 646 0 3 22
0 32 24 34
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
3189 0 0
2
42661.1 0
0
5 4081~
219 1605 591 0 3 22
0 36 35 24
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
8460 0 0
2
42661.1 0
0
9 4-In AND~
219 1490 1070 0 5 22
0 40 39 38 37 144
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 HLT
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 8 0
1 U
5179 0 0
2
42661.1 0
0
9 4-In AND~
219 1488 1018 0 5 22
0 44 43 41 42 12
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 OUT
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 8 0
1 U
3593 0 0
2
42661.1 0
0
9 4-In AND~
219 1489 962 0 5 22
0 44 43 41 37 35
0
0 0 624 0
6 74LS21
-21 -28 21 -20
2 JZ
-8 -28 6 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 18
65 0 0 0 2 2 7 0
1 U
3928 0 0
2
42661.1 0
0
9 4-In AND~
219 1485 910 0 5 22
0 44 43 38 42 25
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 JMP
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
363 0 0
2
42661.1 0
0
9 4-In AND~
219 1483 859 0 5 22
0 44 43 38 37 18
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 MOV
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 6 0
1 U
8132 0 0
2
42661.1 0
0
9 4-In AND~
219 1479 802 0 5 22
0 44 39 41 42 19
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 AND
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 6 0
1 U
65 0 0
2
42661.1 0
0
9 4-In AND~
219 1478 746 0 5 22
0 44 39 41 37 20
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 SUB
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
6609 0 0
2
42661.1 0
0
9 4-In AND~
219 1472 685 0 5 22
0 44 39 38 42 21
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 ADD
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
8995 0 0
2
42661.1 0
0
9 4-In AND~
219 1467 633 0 5 22
0 44 39 38 37 31
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 LOAD
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
3918 0 0
2
42661.1 0
0
7 Ground~
168 113 160 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7519 0 0
2
42661 23
0
14 Logic Display~
6 1039 1407 0 1 2
10 95
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
377 0 0
2
42661 24
0
14 Logic Display~
6 968 1390 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8816 0 0
2
42661 25
0
14 Logic Display~
6 982 2319 0 1 2
10 46
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3877 0 0
2
42661 26
0
14 Logic Display~
6 960 2309 0 1 2
10 47
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
926 0 0
2
42661 27
0
14 Logic Display~
6 938 2301 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7262 0 0
2
42661 28
0
14 Logic Display~
6 891 2291 0 1 2
10 49
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5267 0 0
2
42661 29
0
9 Inverter~
13 596 1578 0 2 22
0 58 57
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U10F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
8838 0 0
2
5.89774e-315 5.26354e-315
0
9 Inverter~
13 591 1493 0 2 22
0 50 52
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U10E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
7159 0 0
2
5.89774e-315 5.30499e-315
0
9 Inverter~
13 600 1551 0 2 22
0 56 55
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U10D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
5812 0 0
2
5.89774e-315 5.32571e-315
0
9 Inverter~
13 609 1532 0 2 22
0 54 53
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U10C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
331 0 0
2
5.89774e-315 5.34643e-315
0
7 Pulser~
4 1797 228 0 11 12
0 61 60 59 145 0 0 10 10 -1
7 1
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 1 0 0
1 V
9604 0 0
2
5.89774e-315 5.3568e-315
0
14 Logic Display~
6 667 1561 0 1 2
10 62
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L102
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7518 0 0
2
42661 30
0
14 Logic Display~
6 843 1497 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L96
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4832 0 0
2
42661 31
0
14 Logic Display~
6 813 1480 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L97
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6798 0 0
2
42661 32
0
14 Logic Display~
6 759 1460 0 1 2
10 64
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L95
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3336 0 0
2
42661 33
0
14 Logic Display~
6 740 1443 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L94
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8370 0 0
2
42661 34
0
14 Logic Display~
6 590 1640 0 1 2
10 66
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L93
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3910 0 0
2
42661 35
0
14 Logic Display~
6 564 1616 0 1 2
10 67
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L92
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
316 0 0
2
42661 36
0
14 Logic Display~
6 535 1597 0 1 2
10 68
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L91
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
536 0 0
2
42661 37
0
14 Logic Display~
6 510 1577 0 1 2
10 69
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L90
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4460 0 0
2
42661 38
0
14 Logic Display~
6 351 1612 0 1 2
10 70
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L89
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3260 0 0
2
42661 39
0
14 Logic Display~
6 323 1583 0 1 2
10 71
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L88
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5156 0 0
2
42661 40
0
14 Logic Display~
6 316 1550 0 1 2
10 72
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L87
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3133 0 0
2
42661 41
0
14 Logic Display~
6 293 1513 0 1 2
10 73
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L86
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
42661 42
0
14 Logic Display~
6 305 1346 0 1 2
10 74
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L85
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3746 0 0
2
5.89774e-315 5.36716e-315
0
14 Logic Display~
6 428 1292 0 1 2
10 75
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L84
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5668 0 0
2
5.89774e-315 5.37752e-315
0
14 Logic Display~
6 407 1284 0 1 2
10 76
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L83
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5368 0 0
2
5.89774e-315 5.38788e-315
0
14 Logic Display~
6 395 1276 0 1 2
10 77
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L82
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8293 0 0
2
5.89774e-315 5.39306e-315
0
14 Logic Display~
6 378 1267 0 1 2
10 78
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L81
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3232 0 0
2
5.89774e-315 5.39824e-315
0
14 Logic Display~
6 528 125 0 1 2
10 79
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L80
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6644 0 0
2
42661 43
0
14 Logic Display~
6 501 115 0 1 2
10 80
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L79
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4978 0 0
2
42661 44
0
14 Logic Display~
6 488 108 0 1 2
10 81
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L78
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9207 0 0
2
42661 45
0
14 Logic Display~
6 475 98 0 1 2
10 82
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L77
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6998 0 0
2
42661 46
0
14 Logic Display~
6 626 2340 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L76
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3175 0 0
2
42661 47
0
14 Logic Display~
6 586 2356 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L75
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3378 0 0
2
42661 48
0
14 Logic Display~
6 546 2375 0 1 2
10 64
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L74
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
922 0 0
2
42661 49
0
14 Logic Display~
6 511 2393 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L73
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6891 0 0
2
42661 50
0
14 Logic Display~
6 247 1218 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L67
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5407 0 0
2
5.89774e-315 5.40342e-315
0
14 Logic Display~
6 227 1213 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L66
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7349 0 0
2
5.89774e-315 5.4086e-315
0
14 Logic Display~
6 215 1208 0 1 2
10 64
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L65
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3919 0 0
2
5.89774e-315 5.41378e-315
0
14 Logic Display~
6 200 1196 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L64
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9747 0 0
2
5.89774e-315 5.41896e-315
0
14 Logic Display~
6 2273 1504 0 1 2
10 74
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L57
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5310 0 0
2
5.89774e-315 5.42414e-315
0
5 4049~
219 2398 1428 0 2 22
0 8 83
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U15E
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 12 0
1 U
4318 0 0
2
42661 51
0
5 4049~
219 2346 1445 0 2 22
0 11 84
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U15D
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 12 0
1 U
3917 0 0
2
42661 52
0
5 4049~
219 2197 1445 0 2 22
0 14 85
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U15C
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 12 0
1 U
7930 0 0
2
42661 53
0
5 4049~
219 2114 1444 0 2 22
0 22 86
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U15B
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 12 0
1 U
6128 0 0
2
42661 54
0
5 4049~
219 2044 1445 0 2 22
0 28 87
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U15A
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 12 0
1 U
7346 0 0
2
42661 55
0
5 4049~
219 1971 1445 0 2 22
0 29 3
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12F
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
8577 0 0
2
42661 56
0
5 4049~
219 1914 1446 0 2 22
0 33 88
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12E
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3372 0 0
2
42661 57
0
14 Logic Display~
6 2349 1486 0 1 2
10 84
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L63
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3741 0 0
2
42661 58
0
14 Logic Display~
6 2421 1485 0 1 2
10 83
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L62
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5813 0 0
2
42661 59
0
14 Logic Display~
6 2574 1481 0 1 2
10 4
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L61
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3213 0 0
2
42661 60
0
14 Logic Display~
6 2502 1482 0 1 2
10 17
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L60
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3694 0 0
2
42661 61
0
14 Logic Display~
6 2047 1492 0 1 2
10 87
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L59
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4327 0 0
2
42661 62
0
14 Logic Display~
6 2119 1498 0 1 2
10 86
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L58
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8800 0 0
2
42661 63
0
14 Logic Display~
6 2200 1488 0 1 2
10 85
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L56
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3406 0 0
2
42661 64
0
14 Logic Display~
6 1902 1493 0 1 2
10 88
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L55
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6455 0 0
2
42661 65
0
14 Logic Display~
6 1974 1492 0 1 2
10 3
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L54
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9319 0 0
2
42661 66
0
14 Logic Display~
6 1821 1496 0 1 2
10 27
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L53
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3172 0 0
2
42661 67
0
14 Logic Display~
6 1749 1497 0 1 2
10 28
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L52
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
38 0 0
2
42661 68
0
5 4049~
219 1339 133 0 2 22
0 42 37
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12D
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
376 0 0
2
42661 69
0
5 4049~
219 1302 130 0 2 22
0 41 38
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12C
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
6666 0 0
2
42661 70
0
5 4049~
219 1259 132 0 2 22
0 43 39
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12B
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
9365 0 0
2
42661 71
0
5 4049~
219 1212 129 0 2 22
0 40 44
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12A
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3251 0 0
2
42661 72
0
14 Logic Display~
6 1210 2276 0 1 2
10 44
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5481 0 0
2
42661 73
0
14 Logic Display~
6 1261 2275 0 1 2
10 39
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L41
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7788 0 0
2
42661 74
0
14 Logic Display~
6 1314 2272 0 1 2
10 38
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L42
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3273 0 0
2
42661 75
0
14 Logic Display~
6 1367 2276 0 1 2
10 37
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L39
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3761 0 0
2
42661 76
0
14 Logic Display~
6 2685 548 0 1 2
10 30
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L38
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
42661 77
0
14 Logic Display~
6 2681 487 0 1 2
10 28
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L37
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4244 0 0
2
42661 78
0
14 Logic Display~
6 2680 417 0 1 2
10 13
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L36
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5225 0 0
2
42661 79
0
14 Logic Display~
6 2677 360 0 1 2
10 32
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L35
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
768 0 0
2
42661 80
0
7 74LS107
112 2398 235 0 12 25
0 30 92 59 89 94 32 59 89 28
91 92 30
0
0 0 4848 0
7 74LS107
-24 -51 25 -43
2 U6
-8 -52 6 -44
0
15 DVCC=14;DGND=7;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 4 12 13 8 11 9 10 3
2 5 6 1 4 12 13 8 11 9
10 3 2 5 6 0
65 0 0 0 1 0 0 0
1 U
5735 0 0
2
42661 81
0
7 74LS107
112 2179 243 0 12 25
0 13 93 59 89 28 91 59 89 32
94 13 93
0
0 0 4848 0
7 74LS107
-24 -51 25 -43
2 U1
-8 -52 6 -44
0
15 DVCC=14;DGND=7;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 4 12 13 8 11 9 10 3
2 5 6 1 4 12 13 8 11 9
10 3 2 5 6 0
65 0 0 0 1 0 0 0
1 U
5881 0 0
2
42661 82
0
7 74LS173
129 574 2300 0 14 29
0 2 84 84 90 65 64 45 63 2
2 49 48 47 46
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3275 0 0
2
42661 83
0
7 Ground~
168 528 2128 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4203 0 0
2
42661 84
0
9 Inverter~
13 675 2128 0 2 22
0 96 69
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U10B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3440 0 0
2
42661 85
0
9 Inverter~
13 673 2087 0 2 22
0 97 68
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U10A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
9102 0 0
2
42661 86
0
9 Inverter~
13 633 2021 0 2 22
0 98 66
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
5586 0 0
2
42661 87
0
9 Inverter~
13 622 1975 0 2 22
0 99 67
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
525 0 0
2
42661 88
0
7 74LS173
129 408 2210 0 14 29
0 2 2 2 90 112 111 110 109 2
2 105 106 107 108
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6206 0 0
2
42661 89
0
7 74LS157
122 569 2047 0 14 29
0 100 108 104 107 103 106 102 105 101
2 99 98 97 96
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3418 0 0
2
42661 90
0
7 74LS126
116 568 1772 0 12 25
0 17 101 17 102 17 103 17 104 65
64 45 63
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U7
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
9312 0 0
2
42661 91
0
7 Ground~
168 364 1908 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7419 0 0
2
42661 92
0
7 74LS173
129 428 1772 0 14 29
0 2 2 2 90 116 115 114 113 2
2 101 102 103 104
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
472 0 0
2
42661 93
0
7 74LS126
116 707 1478 0 12 25
0 62 51 62 53 62 55 62 57 65
64 45 63
0
0 0 4848 0
7 74LS126
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
4714 0 0
2
42661 94
0
9 Inverter~
13 241 1628 0 2 22
0 75 70
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9386 0 0
2
42661 95
0
9 Inverter~
13 241 1599 0 2 22
0 76 71
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
7610 0 0
2
42661 96
0
9 Inverter~
13 242 1567 0 2 22
0 77 72
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3482 0 0
2
42661 97
0
9 Inverter~
13 243 1531 0 2 22
0 78 73
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3608 0 0
2
42661 98
0
7 74LS181
132 518 1474 0 22 45
0 122 121 120 119 73 72 71 70 69
68 66 67 118 117 95 36 146 147 50
54 56 58
0
0 0 4848 0
7 74LS181
-24 -69 25 -61
2 U3
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
6397 0 0
2
42661 99
0
7 Ground~
168 168 1248 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3967 0 0
2
42661 100
0
7 74LS126
116 533 1274 0 12 25
0 74 78 74 77 74 76 74 75 65
64 45 63
0
0 0 4848 0
7 74LS126
-24 -51 25 -43
3 ACC
-10 -52 11 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
8621 0 0
2
42661 101
0
7 74LS173
129 310 1276 0 14 29
0 2 85 85 90 65 64 45 63 2
2 78 77 76 75
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
3 ACC
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
8901 0 0
2
42661 102
0
14 Logic Display~
6 666 1023 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L28
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7385 0 0
2
42661 103
0
14 Logic Display~
6 646 1013 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L27
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6519 0 0
2
42661 104
0
14 Logic Display~
6 625 1005 0 1 2
10 64
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L26
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
552 0 0
2
42661 105
0
14 Logic Display~
6 597 997 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L25
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
42661 106
0
7 Ground~
168 388 998 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8715 0 0
2
42661 107
0
14 Logic Display~
6 419 1129 0 1 2
10 42
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L24
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9763 0 0
2
42661 108
0
14 Logic Display~
6 374 1124 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L23
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8443 0 0
2
42661 109
0
14 Logic Display~
6 337 1126 0 1 2
10 43
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L22
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3719 0 0
2
42661 110
0
14 Logic Display~
6 302 1127 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L21
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8671 0 0
2
42661 111
0
7 74LS173
129 515 1004 0 14 29
0 2 87 87 90 65 64 45 63 86
86 65 64 45 63
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
2 IR
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
42661 112
0
7 74LS173
129 321 1004 0 14 29
0 2 87 87 90 126 125 124 123 2
2 40 43 41 42
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
2 IR
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
49 0 0
2
42661 113
0
2 +V
167 597 758 0 1 3
0 128
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6536 0 0
2
42661 114
0
14 Logic Display~
6 850 844 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L20
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3931 0 0
2
42661 115
0
14 Logic Display~
6 822 833 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4390 0 0
2
42661 116
0
14 Logic Display~
6 790 826 0 1 2
10 64
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3242 0 0
2
42661 117
0
14 Logic Display~
6 763 817 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6760 0 0
2
42661 118
0
14 Logic Display~
6 733 807 0 1 2
10 123
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5760 0 0
2
42661 119
0
14 Logic Display~
6 712 799 0 1 2
10 124
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3781 0 0
2
42661 120
0
14 Logic Display~
6 681 788 0 1 2
10 125
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8545 0 0
2
42661 121
0
14 Logic Display~
6 639 779 0 1 2
10 126
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9739 0 0
2
42661 122
0
7 Ground~
168 370 778 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
388 0 0
2
42661 0
0
6 1K RAM
79 487 815 0 20 41
0 129 129 129 129 129 129 130 131 127
132 126 125 124 123 65 64 45 63 3
128
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U2
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 1 0 0 0
1 U
4595 0 0
2
42661 1
0
14 Logic Display~
6 604 566 0 1 2
10 130
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3173 0 0
2
42661 2
0
14 Logic Display~
6 583 564 0 1 2
10 131
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9261 0 0
2
42661 3
0
14 Logic Display~
6 556 568 0 1 2
10 127
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3494 0 0
2
42661 4
0
14 Logic Display~
6 532 570 0 1 2
10 132
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9101 0 0
2
42661 5
0
7 Ground~
168 430 684 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
358 0 0
2
42661 6
0
7 74LS157
122 488 605 0 14 29
0 137 136 141 135 140 134 139 133 138
2 132 127 131 130
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3726 0 0
2
42661 7
0
7 74LS173
129 495 397 0 14 29
0 2 88 88 90 65 64 45 63 2
2 138 139 140 141
0
0 0 4848 0
7 74LS173
-24 -51 25 -43
3 MAR
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
999 0 0
2
42661 8
0
7 Ground~
168 323 183 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8787 0 0
2
5.89774e-315 5.42933e-315
0
7 74LS126
116 588 106 0 12 25
0 27 82 27 81 27 80 27 79 65
64 45 63
0
0 0 4848 0
7 74LS126
-24 -51 25 -43
2 PC
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3348 0 0
2
5.89774e-315 5.43192e-315
0
7 74LS193
137 426 106 0 14 29
0 90 28 83 2 65 64 45 63 148
149 82 81 80 79
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 PC
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3395 0 0
2
5.89774e-315 5.43451e-315
0
7 Pulser~
4 176 72 0 11 12
0 143 142 90 150 0 0 10 10 -1
7 1
0
0 0 4656 0
0
3 V20
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 1 0 0
1 V
7740 0 0
2
5.89774e-315 5.4371e-315
0
414
1 4 4 0 0 4224 0 106 25 0 0 4
2574 1467
2574 868
2553 868
2553 852
0 3 5 0 0 4224 0 0 25 15 0 3
2177 793
2544 793
2544 806
0 2 6 0 0 4224 0 0 25 16 0 3
2186 739
2553 739
2553 807
0 1 7 0 0 4224 0 0 25 17 0 3
2162 683
2562 683
2562 806
3 1 8 0 0 4224 0 26 97 0 0 3
2379 1050
2379 1410
2401 1410
3 1 9 0 0 4224 0 36 26 0 0 3
2099 909
2388 909
2388 1004
0 2 10 0 0 4224 0 0 26 27 0 3
2088 976
2370 976
2370 1004
0 3 11 0 0 4224 0 0 27 156 0 2
2274 1423
2274 828
5 2 12 0 0 4224 0 46 27 0 0 3
1509 1018
2229 1018
2229 837
1 0 13 0 0 4096 0 27 0 0 195 4
2229 819
2229 444
2244 444
2244 429
1 3 14 0 0 12416 0 99 28 0 0 4
2200 1427
2200 1412
2210 1412
2210 1033
5 1 15 0 0 4224 0 29 28 0 0 3
2182 961
2219 961
2219 987
0 2 16 0 0 8320 0 0 28 42 0 3
1966 650
2201 650
2201 987
4 3 17 0 0 4096 0 29 30 0 0 3
2168 911
2168 851
2163 851
3 3 5 0 0 0 0 31 29 0 0 3
2161 793
2177 793
2177 911
2 3 6 0 0 0 0 29 32 0 0 4
2186 911
2186 739
2172 739
2172 746
1 3 7 0 0 0 0 29 33 0 0 4
2195 911
2195 893
2162 893
2162 679
5 2 18 0 0 12416 0 49 30 0 0 4
1504 859
1519 859
1519 860
2118 860
0 1 13 0 0 0 0 0 30 21 0 3
1775 784
1775 842
2118 842
5 2 19 0 0 4224 0 50 31 0 0 2
1500 802
2116 802
0 1 13 0 0 0 0 0 31 23 0 3
1775 737
1775 784
2116 784
5 2 20 0 0 12416 0 51 32 0 0 5
1499 746
1605 746
1605 759
2127 759
2127 755
0 1 13 0 0 0 0 0 32 49 0 3
1775 591
1775 737
2127 737
1 0 13 0 0 0 0 33 0 0 195 4
2117 670
2117 444
2145 444
2145 429
5 2 21 0 0 12416 0 52 33 0 0 5
1493 685
1604 685
1604 719
2117 719
2117 688
1 4 22 0 0 8320 0 100 34 0 0 3
2117 1426
2097 1426
2097 1041
3 3 10 0 0 0 0 34 35 0 0 3
2088 995
2088 976
2076 976
1 3 23 0 0 4224 0 34 40 0 0 3
2106 995
2106 602
1851 602
2 3 9 0 0 0 0 34 36 0 0 3
2097 996
2097 909
2099 909
0 2 24 0 0 8320 0 0 35 56 0 3
1626 655
1626 985
2031 985
0 1 13 0 0 0 0 0 35 33 0 5
2067 745
2067 744
2021 744
2021 967
2031 967
0 2 25 0 0 16512 0 0 36 54 0 5
1649 910
1649 917
1707 917
1707 918
2054 918
1 0 13 0 0 8192 0 36 0 0 195 3
2054 900
2067 900
2067 429
0 4 26 0 0 4224 0 0 39 40 0 3
1755 696
1866 696
1866 633
0 0 27 0 0 4096 0 0 0 39 51 2
1821 1470
1791 1470
0 1 28 0 0 8192 0 0 101 41 0 3
1988 619
2047 619
2047 1427
1 3 29 0 0 4224 0 102 37 0 0 3
1974 1427
1974 752
1957 752
0 2 30 0 0 4096 0 0 41 193 0 3
1740 560
1740 667
1764 667
1 4 27 0 0 4096 0 113 41 0 0 3
1821 1482
1821 667
1809 667
3 3 26 0 0 0 0 42 41 0 0 4
1714 696
1758 696
1758 676
1763 676
0 2 28 0 0 0 0 0 37 194 0 4
1988 499
1988 687
1948 687
1948 706
1 3 16 0 0 0 0 37 38 0 0 3
1966 706
1966 649
1969 649
0 2 31 0 0 8192 0 0 38 50 0 3
1793 611
1793 658
1924 658
0 1 32 0 0 4096 0 0 38 196 0 3
1922 372
1922 640
1924 640
1 5 33 0 0 4224 0 103 39 0 0 4
1917 1428
1917 672
1916 672
1916 619
0 1 30 0 0 0 0 0 39 193 0 3
1861 560
1861 606
1866 606
0 3 34 0 0 8320 0 0 39 53 0 3
1758 646
1758 624
1866 624
3 2 23 0 0 0 0 40 39 0 0 4
1851 602
1851 614
1866 614
1866 615
0 1 13 0 0 0 0 0 40 195 0 3
1775 429
1775 593
1806 593
2 5 31 0 0 4224 0 40 53 0 0 4
1806 611
1499 611
1499 633
1488 633
0 0 27 0 0 0 0 0 0 0 406 2
1817 1470
1791 1470
0 2 28 0 0 24704 0 0 180 61 0 8
1749 1479
1742 1479
1742 2184
1928 2184
1928 2644
6 2644
6 88
394 88
3 1 34 0 0 0 0 43 41 0 0 4
1707 646
1758 646
1758 658
1763 658
5 2 25 0 0 0 0 48 42 0 0 4
1506 910
1649 910
1649 705
1669 705
0 1 32 0 0 0 0 0 42 57 0 4
1662 600
1650 600
1650 687
1669 687
3 2 24 0 0 0 0 44 43 0 0 3
1626 591
1626 655
1662 655
0 1 32 0 0 0 0 0 43 196 0 4
1864 372
1864 393
1662 393
1662 637
5 2 35 0 0 8320 0 47 44 0 0 4
1510 962
1579 962
1579 600
1581 600
0 0 36 0 0 4096 0 0 0 198 60 2
1019 167
1019 411
0 1 36 0 0 4224 0 0 44 100 0 5
1019 1327
1019 411
1567 411
1567 582
1581 582
1 0 28 0 0 0 0 114 0 0 194 2
1749 1483
1749 499
4 0 37 0 0 4096 0 45 0 0 165 2
1466 1084
1367 1084
3 0 38 0 0 4096 0 45 0 0 166 2
1466 1075
1305 1075
2 0 39 0 0 4096 0 45 0 0 167 2
1466 1066
1262 1066
1 0 40 0 0 4096 0 45 0 0 199 2
1466 1057
1193 1057
4 0 37 0 0 0 0 47 0 0 165 2
1465 976
1367 976
3 0 41 0 0 4096 0 47 0 0 201 2
1465 967
1289 967
4 0 42 0 0 4096 0 46 0 0 202 2
1464 1032
1347 1032
3 0 41 0 0 0 0 46 0 0 201 2
1464 1023
1289 1023
2 0 43 0 0 4096 0 46 0 0 200 2
1464 1014
1244 1014
1 0 44 0 0 4096 0 46 0 0 168 2
1464 1005
1215 1005
2 0 43 0 0 4096 0 47 0 0 200 2
1465 958
1244 958
1 0 44 0 0 4096 0 47 0 0 168 2
1465 949
1215 949
4 0 42 0 0 0 0 48 0 0 202 2
1461 924
1347 924
3 0 38 0 0 0 0 48 0 0 166 2
1461 915
1305 915
2 0 43 0 0 0 0 48 0 0 200 2
1461 906
1244 906
1 0 44 0 0 0 0 48 0 0 168 2
1461 897
1215 897
4 0 37 0 0 0 0 49 0 0 165 2
1459 873
1367 873
3 0 38 0 0 0 0 49 0 0 166 2
1459 864
1305 864
2 0 43 0 0 0 0 49 0 0 200 2
1459 855
1244 855
1 0 44 0 0 0 0 49 0 0 168 2
1459 846
1215 846
4 0 42 0 0 0 0 50 0 0 202 2
1455 816
1347 816
3 0 41 0 0 0 0 50 0 0 201 2
1455 807
1289 807
2 0 39 0 0 0 0 50 0 0 167 2
1455 798
1262 798
1 0 44 0 0 0 0 50 0 0 168 2
1455 789
1215 789
4 0 37 0 0 0 0 51 0 0 165 2
1454 760
1367 760
3 0 41 0 0 0 0 51 0 0 201 2
1454 751
1289 751
2 0 39 0 0 0 0 51 0 0 167 2
1454 742
1262 742
1 0 44 0 0 0 0 51 0 0 168 2
1454 733
1215 733
4 0 42 0 0 0 0 52 0 0 202 2
1448 699
1347 699
3 0 38 0 0 0 0 52 0 0 166 2
1448 690
1305 690
2 0 39 0 0 0 0 52 0 0 167 2
1448 681
1262 681
1 0 44 0 0 0 0 52 0 0 168 2
1448 672
1215 672
4 0 37 0 0 0 0 53 0 0 165 2
1443 647
1367 647
3 0 38 0 0 0 0 53 0 0 166 2
1443 638
1305 638
2 0 39 0 0 0 0 53 0 0 167 2
1443 629
1262 629
1 0 44 0 0 0 0 53 0 0 168 2
1443 620
1215 620
0 0 45 0 0 4096 0 0 0 269 309 2
829 1299
829 1187
0 1 2 0 0 4096 0 0 54 132 0 2
114 141
113 154
16 0 36 0 0 128 0 145 0 0 0 9
550 1474
610 1474
610 1450
594 1450
594 1443
621 1443
621 1407
1019 1407
1019 1324
1 0 36 0 0 0 0 56 0 0 100 2
968 1408
968 1407
1 0 46 0 0 4096 0 57 0 0 206 2
982 2337
982 2336
1 0 47 0 0 0 0 58 0 0 205 2
960 2327
960 2327
1 0 48 0 0 4096 0 59 0 0 204 2
938 2319
938 2318
1 0 49 0 0 0 0 60 0 0 203 2
891 2309
891 2309
19 1 50 0 0 4224 0 145 62 0 0 3
556 1501
576 1501
576 1493
2 0 51 0 0 4224 0 140 0 0 0 2
675 1460
628 1460
2 0 52 0 0 8320 0 62 0 0 0 3
612 1493
628 1493
628 1460
2 4 53 0 0 8320 0 64 140 0 0 4
630 1532
631 1532
631 1478
675 1478
20 1 54 0 0 4224 0 145 64 0 0 3
556 1510
594 1510
594 1532
2 6 55 0 0 8320 0 63 140 0 0 4
621 1551
637 1551
637 1496
675 1496
21 1 56 0 0 8320 0 145 63 0 0 3
556 1519
585 1519
585 1551
2 8 57 0 0 8320 0 61 140 0 0 4
617 1578
645 1578
645 1514
675 1514
22 1 58 0 0 8320 0 145 61 0 0 4
556 1528
562 1528
562 1578
581 1578
0 3 59 0 0 8192 0 0 128 0 0 3
2002 238
2002 234
2141 234
3 1 59 0 0 4096 0 65 0 0 115 3
1821 219
2015 219
2015 234
0 2 60 0 0 4224 0 0 65 0 0 3
1766 232
1766 228
1767 228
1 1 61 0 0 4224 0 65 1 0 0 4
1773 219
1739 219
1739 227
1726 227
1 0 62 0 0 4096 0 66 0 0 274 2
667 1579
668 1579
1 0 63 0 0 4096 0 67 0 0 270 2
843 1515
843 1514
1 0 45 0 0 0 0 68 0 0 269 2
813 1498
813 1496
1 0 64 0 0 0 0 69 0 0 268 2
759 1478
759 1478
1 0 65 0 0 4096 0 70 0 0 267 2
740 1461
740 1460
1 0 66 0 0 4096 0 71 0 0 223 2
590 1658
590 1657
1 0 67 0 0 0 0 72 0 0 224 2
564 1634
564 1634
1 0 68 0 0 4096 0 73 0 0 222 2
535 1615
535 1613
1 0 69 0 0 4096 0 74 0 0 221 2
510 1595
510 1593
1 0 70 0 0 4096 0 75 0 0 275 2
351 1630
351 1628
1 0 71 0 0 4096 0 76 0 0 276 2
323 1601
323 1599
1 0 72 0 0 4096 0 77 0 0 277 2
316 1568
316 1567
1 0 73 0 0 0 0 78 0 0 278 2
293 1531
293 1531
0 4 2 0 0 12288 0 0 180 0 0 4
114 141
174 141
174 106
394 106
1 0 74 0 0 4096 0 79 0 0 296 2
305 1364
305 1365
1 0 75 0 0 0 0 80 0 0 300 2
428 1310
428 1310
1 0 76 0 0 4096 0 81 0 0 299 2
407 1302
407 1303
1 0 77 0 0 0 0 82 0 0 298 2
395 1294
395 1294
1 0 78 0 0 0 0 83 0 0 297 2
378 1285
378 1285
1 0 79 0 0 4096 0 84 0 0 411 2
528 143
528 142
1 0 80 0 0 0 0 85 0 0 410 2
501 133
501 133
1 0 81 0 0 4096 0 86 0 0 409 2
488 126
488 124
1 0 82 0 0 4096 0 87 0 0 408 2
475 116
475 115
1 0 63 0 0 4096 0 88 0 0 216 2
626 2358
626 2356
1 0 45 0 0 0 0 89 0 0 215 2
586 2374
586 2372
1 0 64 0 0 4096 0 90 0 0 214 2
546 2393
546 2391
1 0 65 0 0 0 0 91 0 0 213 2
511 2411
511 2410
0 0 64 0 0 4096 0 0 0 0 291 3
659 1254
659 1274
656 1274
1 0 63 0 0 0 0 92 0 0 310 2
247 1236
247 1236
1 0 45 0 0 0 0 93 0 0 309 2
227 1231
228 1231
1 0 64 0 0 0 0 94 0 0 308 2
215 1226
214 1226
1 0 65 0 0 0 0 95 0 0 307 2
200 1214
200 1214
0 0 17 0 0 12416 0 0 0 252 153 10
193 1972
76 1972
76 2580
1857 2580
1857 2274
1614 2274
1614 1701
2481 1701
2481 1457
2502 1457
0 0 62 0 0 12416 0 0 0 274 0 10
94 1692
64 1692
64 2589
1866 2589
1866 2261
1639 2261
1639 1681
2557 1681
2557 1460
2574 1460
0 1 17 0 0 0 0 0 107 14 0 5
2168 852
2486 852
2486 1426
2502 1426
2502 1468
2 1 83 0 0 8192 0 97 105 0 0 3
2401 1446
2421 1446
2421 1471
2 1 84 0 0 4096 0 98 104 0 0 2
2349 1463
2349 1472
0 1 11 0 0 128 0 0 98 0 0 3
2270 1423
2349 1423
2349 1427
0 1 74 0 0 8192 0 0 96 0 0 3
2270 1423
2273 1423
2273 1490
2 1 85 0 0 4096 0 99 110 0 0 2
2200 1463
2200 1474
2 1 86 0 0 8192 0 100 109 0 0 3
2117 1462
2119 1462
2119 1484
2 1 87 0 0 4096 0 101 108 0 0 2
2047 1463
2047 1478
2 1 3 0 0 4096 0 102 112 0 0 2
1974 1463
1974 1478
2 1 88 0 0 8192 0 103 111 0 0 4
1917 1464
1917 1470
1902 1470
1902 1479
0 0 42 0 0 0 0 0 0 202 0 5
1347 2303
1335 2303
1335 2313
1341 2313
1341 2341
0 0 41 0 0 0 0 0 0 201 0 5
1289 2299
1291 2299
1291 2323
1289 2323
1289 2345
1 2 37 0 0 4224 0 122 115 0 0 3
1367 2262
1367 151
1342 151
2 1 38 0 0 4224 0 116 121 0 0 3
1305 148
1305 2258
1314 2258
1 2 39 0 0 8320 0 120 117 0 0 3
1261 2261
1262 2261
1262 150
2 1 44 0 0 4224 0 118 119 0 0 3
1215 147
1215 2262
1210 2262
1 0 42 0 0 0 0 115 0 0 202 3
1342 115
1342 104
1347 104
1 0 41 0 0 0 0 116 0 0 201 3
1305 112
1305 103
1289 103
1 0 43 0 0 0 0 117 0 0 200 3
1262 114
1262 98
1244 98
1 0 40 0 0 0 0 118 0 0 199 3
1215 111
1215 100
1193 100
0 7 59 0 0 0 0 0 127 174 0 3
2341 225
2341 262
2360 262
0 3 59 0 0 8320 0 0 127 175 0 5
2071 234
2071 183
2341 183
2341 226
2360 226
0 7 59 0 0 0 0 0 128 115 0 3
2071 234
2071 270
2141 270
8 0 89 0 0 4096 0 127 0 0 177 2
2360 271
2311 271
0 4 89 0 0 4224 0 0 127 179 0 4
2028 295
2311 295
2311 235
2360 235
8 0 89 0 0 0 0 128 0 0 179 2
2141 279
2028 279
4 1 89 0 0 0 0 128 3 0 0 4
2141 243
2028 243
2028 296
1798 296
0 0 90 0 0 4224 0 0 0 0 412 3
1716 306
226 306
226 63
6 10 91 0 0 12416 0 128 127 0 0 6
2147 261
2096 261
2096 157
2480 157
2480 226
2436 226
5 0 28 0 0 0 0 128 0 0 184 5
2147 252
2108 252
2108 169
2490 169
2490 217
0 0 30 0 0 4096 0 0 0 185 193 2
2498 262
2498 560
9 0 28 0 0 0 0 127 0 0 194 3
2430 217
2490 217
2490 499
12 1 30 0 0 0 0 127 127 0 0 6
2436 262
2501 262
2501 67
2319 67
2319 208
2366 208
11 2 92 0 0 12416 0 127 127 0 0 6
2430 253
2509 253
2509 59
2311 59
2311 217
2366 217
0 0 13 0 0 0 0 0 0 189 195 2
2229 308
2229 429
12 2 93 0 0 8320 0 128 128 0 0 5
2217 270
2217 300
2130 300
2130 225
2147 225
11 1 13 0 0 0 0 128 128 0 0 6
2211 261
2229 261
2229 309
2121 309
2121 216
2147 216
5 10 94 0 0 4224 0 127 128 0 0 3
2366 244
2217 244
2217 234
6 0 32 0 0 0 0 127 0 0 192 2
2366 253
2247 253
9 0 32 0 0 0 0 128 0 0 196 3
2211 225
2247 225
2247 372
0 1 30 0 0 4224 0 0 123 0 0 4
1733 560
2662 560
2662 552
2669 552
0 1 28 0 0 128 0 0 124 0 0 4
1729 499
2658 499
2658 491
2665 491
0 1 13 0 0 4224 0 0 125 0 0 4
1728 429
2657 429
2657 421
2664 421
0 1 32 0 0 4224 0 0 126 0 0 4
1725 372
2654 372
2654 364
2661 364
1 15 95 0 0 8320 0 55 145 0 0 5
1039 1425
1040 1423
599 1423
599 1465
550 1465
0 1 36 0 0 128 0 0 2 0 0 4
1019 65
1019 167
1148 167
1148 204
1 0 40 0 0 20608 0 157 0 0 0 12
302 1145
302 1154
1110 1154
1110 69
1193 69
1193 2289
1182 2289
1182 2303
1171 2303
1171 2323
1169 2323
1169 2344
1 0 43 0 0 20608 0 156 0 0 0 11
337 1144
337 1150
1096 1150
1096 58
1244 58
1244 2302
1233 2302
1233 2318
1232 2318
1232 2347
1229 2347
0 0 41 0 0 16512 0 0 0 331 0 6
360 1097
1082 1097
1082 41
1289 41
1289 2299
1286 2299
0 0 42 0 0 24704 0 0 0 332 163 8
403 1092
1064 1092
1064 16
1366 16
1366 77
1347 77
1347 2303
1335 2303
0 11 49 0 0 4224 0 0 129 0 0 2
919 2309
606 2309
0 12 48 0 0 4224 0 0 129 0 0 2
947 2318
606 2318
0 13 47 0 0 4224 0 0 129 0 0 2
968 2327
606 2327
0 14 46 0 0 4224 0 0 129 0 0 2
993 2336
606 2336
0 4 90 0 0 0 0 0 129 217 0 3
364 2210
364 2300
542 2300
0 10 2 0 0 0 0 0 129 210 0 4
542 2174
635 2174
635 2282
612 2282
9 0 2 0 0 0 0 129 0 0 210 3
612 2273
612 2187
542 2187
0 1 2 0 0 0 0 0 129 220 0 3
531 2112
542 2112
542 2273
2 0 84 0 0 4096 0 129 0 0 212 3
536 2282
523 2282
523 2291
3 1 84 0 0 20608 0 129 104 0 0 14
536 2291
355 2291
355 2388
109 2388
109 2569
1843 2569
1843 2289
1600 2289
1600 1719
2350 1719
2350 1541
2323 1541
2323 1472
2349 1472
0 5 65 0 0 4224 0 0 129 245 0 5
773 1752
773 2410
496 2410
496 2309
542 2309
0 6 64 0 0 4224 0 0 129 246 0 5
801 1769
801 2391
519 2391
519 2318
542 2318
0 7 45 0 0 4096 0 0 129 247 0 5
829 1790
829 2372
531 2372
531 2327
542 2327
0 8 63 0 0 4096 0 0 129 248 0 4
852 1808
852 2356
542 2356
542 2336
0 4 90 0 0 0 0 0 135 257 0 5
328 1728
328 2146
356 2146
356 2210
376 2210
2 0 2 0 0 0 0 135 0 0 244 2
370 2192
370 2183
0 3 2 0 0 0 0 0 135 244 0 3
363 2183
363 2201
370 2201
10 1 2 0 0 0 0 136 130 0 0 4
531 2092
531 2113
528 2113
528 2122
2 9 69 0 0 8320 0 131 145 0 0 6
696 2128
722 2128
722 1593
427 1593
427 1501
480 1501
2 10 68 0 0 8320 0 132 145 0 0 6
694 2087
704 2087
704 1613
443 1613
443 1510
480 1510
2 11 66 0 0 8320 0 133 145 0 0 6
654 2021
656 2021
656 1657
452 1657
452 1519
480 1519
2 12 67 0 0 4224 0 134 145 0 0 5
643 1975
643 1634
481 1634
481 1528
480 1528
1 14 96 0 0 4224 0 131 136 0 0 4
660 2128
615 2128
615 2083
601 2083
1 13 97 0 0 12416 0 132 136 0 0 4
658 2087
637 2087
637 2065
601 2065
1 12 98 0 0 4224 0 133 136 0 0 3
618 2021
618 2047
601 2047
11 1 99 0 0 8320 0 136 134 0 0 3
601 2029
607 2029
607 1975
1 1 100 0 0 12416 0 4 136 0 0 4
217 2033
306 2033
306 2011
537 2011
0 9 101 0 0 4224 0 0 136 253 0 3
513 1754
513 2083
537 2083
0 7 102 0 0 4224 0 0 136 254 0 3
502 1772
502 2065
537 2065
0 5 103 0 0 4224 0 0 136 255 0 3
495 1799
495 2047
537 2047
0 3 104 0 0 4224 0 0 136 256 0 3
484 1808
484 2029
537 2029
11 8 105 0 0 8320 0 135 136 0 0 4
440 2219
466 2219
466 2074
537 2074
12 6 106 0 0 8320 0 135 136 0 0 4
440 2228
470 2228
470 2056
537 2056
13 4 107 0 0 8320 0 135 136 0 0 4
440 2237
481 2237
481 2038
537 2038
14 2 108 0 0 8320 0 135 136 0 0 4
440 2246
491 2246
491 2020
537 2020
1 8 109 0 0 12416 0 5 135 0 0 4
214 2293
238 2293
238 2246
376 2246
1 7 110 0 0 12416 0 6 135 0 0 4
216 2247
226 2247
226 2237
376 2237
1 6 111 0 0 12416 0 7 135 0 0 4
216 2203
235 2203
235 2228
376 2228
1 5 112 0 0 12416 0 8 135 0 0 4
216 2158
278 2158
278 2219
376 2219
9 0 2 0 0 0 0 135 0 0 243 2
446 2183
453 2183
0 10 2 0 0 0 0 0 135 244 0 5
393 2119
393 2149
453 2149
453 2192
446 2192
0 1 2 0 0 8320 0 0 135 262 0 6
364 1877
393 1877
393 2120
360 2120
360 2183
376 2183
0 9 65 0 0 0 0 0 137 267 0 3
773 1460
773 1754
600 1754
0 10 64 0 0 0 0 0 137 268 0 3
801 1478
801 1772
600 1772
0 11 45 0 0 0 0 0 137 269 0 3
829 1493
829 1790
600 1790
0 12 63 0 0 0 0 0 137 270 0 3
852 1514
852 1808
600 1808
7 0 17 0 0 0 0 137 0 0 252 2
536 1799
522 1799
5 0 17 0 0 0 0 137 0 0 252 2
536 1781
522 1781
3 0 17 0 0 0 0 137 0 0 252 2
536 1763
522 1763
0 1 17 0 0 0 0 0 137 0 0 4
185 1972
522 1972
522 1745
536 1745
11 2 101 0 0 0 0 139 137 0 0 4
460 1781
491 1781
491 1754
536 1754
12 4 102 0 0 0 0 139 137 0 0 4
460 1790
478 1790
478 1772
536 1772
13 6 103 0 0 0 0 139 137 0 0 4
460 1799
496 1799
496 1790
536 1790
14 8 104 0 0 0 0 139 137 0 0 2
460 1808
536 1808
0 4 90 0 0 0 0 0 139 306 0 6
102 1276
130 1276
130 1728
334 1728
334 1772
396 1772
10 9 2 0 0 0 0 139 139 0 0 5
466 1754
480 1754
480 1738
466 1738
466 1745
0 9 2 0 0 0 0 0 139 260 0 4
365 1745
365 1703
466 1703
466 1745
1 0 2 0 0 0 0 139 0 0 262 3
396 1745
364 1745
364 1754
3 0 2 0 0 0 0 139 0 0 262 2
390 1763
364 1763
2 1 2 0 0 0 0 139 138 0 0 3
390 1754
364 1754
364 1902
1 8 113 0 0 4224 0 9 139 0 0 4
223 1888
337 1888
337 1808
396 1808
1 7 114 0 0 4224 0 10 139 0 0 4
222 1850
320 1850
320 1799
396 1799
1 6 115 0 0 12416 0 11 139 0 0 4
223 1813
272 1813
272 1790
396 1790
1 5 116 0 0 12416 0 12 139 0 0 4
222 1772
289 1772
289 1781
396 1781
9 0 65 0 0 0 0 140 0 0 290 3
739 1460
776 1460
776 1234
0 10 64 0 0 0 0 0 140 291 0 3
801 1274
801 1478
739 1478
11 11 45 0 0 0 0 147 140 0 0 6
565 1292
664 1292
664 1299
829 1299
829 1496
739 1496
12 0 63 0 0 0 0 140 0 0 292 3
739 1514
855 1514
855 1310
7 0 62 0 0 0 0 140 0 0 274 2
675 1505
668 1505
5 0 62 0 0 0 0 140 0 0 274 2
675 1487
668 1487
3 0 62 0 0 0 0 140 0 0 274 2
675 1469
668 1469
0 1 62 0 0 0 0 0 140 0 0 4
89 1692
668 1692
668 1451
675 1451
2 8 70 0 0 4224 0 141 145 0 0 4
262 1628
404 1628
404 1492
480 1492
2 7 71 0 0 4224 0 142 145 0 0 4
262 1599
396 1599
396 1483
480 1483
2 6 72 0 0 4224 0 143 145 0 0 4
263 1567
380 1567
380 1474
480 1474
2 5 73 0 0 12416 0 144 145 0 0 4
264 1531
365 1531
365 1465
480 1465
1 0 78 0 0 16512 0 144 0 0 297 5
228 1531
213 1531
213 1514
361 1514
361 1285
1 0 77 0 0 16512 0 143 0 0 298 5
227 1567
199 1567
199 1511
353 1511
353 1294
1 0 76 0 0 16512 0 142 0 0 299 5
226 1599
193 1599
193 1505
347 1505
347 1303
14 0 75 0 0 4096 0 148 0 0 300 2
342 1312
342 1310
1 14 75 0 0 16512 0 141 148 0 0 5
226 1628
182 1628
182 1501
342 1501
342 1312
1 14 117 0 0 8320 0 13 145 0 0 7
210 1416
210 1382
463 1382
463 1372
613 1372
613 1438
550 1438
1 13 118 0 0 4224 0 14 145 0 0 3
208 1389
550 1389
550 1429
1 4 119 0 0 12416 0 15 145 0 0 4
268 1489
287 1489
287 1456
486 1456
3 1 120 0 0 4224 0 145 16 0 0 3
486 1447
268 1447
268 1464
1 2 121 0 0 4224 0 17 145 0 0 3
270 1439
486 1439
486 1438
1 1 122 0 0 4224 0 18 145 0 0 3
270 1414
486 1414
486 1429
0 9 65 0 0 0 0 0 147 307 0 4
776 1159
776 1234
565 1234
565 1256
10 0 64 0 0 0 0 147 0 0 308 3
565 1274
803 1274
803 1177
12 0 63 0 0 0 0 147 0 0 310 3
565 1310
855 1310
855 1207
7 0 74 0 0 0 0 147 0 0 296 2
501 1301
464 1301
5 0 74 0 0 0 0 147 0 0 296 2
501 1283
464 1283
3 0 74 0 0 0 0 147 0 0 296 2
501 1265
464 1265
0 1 74 0 0 32896 0 0 147 157 0 13
2273 1472
2273 1473
2249 1473
2249 1671
1647 1671
1647 2254
1873 2254
1873 2594
56 2594
56 1365
464 1365
464 1247
501 1247
11 2 78 0 0 0 0 148 147 0 0 4
342 1285
407 1285
407 1256
501 1256
12 4 77 0 0 0 0 148 147 0 0 4
342 1294
424 1294
424 1274
501 1274
13 6 76 0 0 0 0 148 147 0 0 4
342 1303
434 1303
434 1292
501 1292
14 8 75 0 0 0 0 148 147 0 0 3
342 1312
342 1310
501 1310
9 0 2 0 0 0 0 148 0 0 302 2
348 1249
363 1249
0 10 2 0 0 0 0 0 148 303 0 5
278 1242
278 1220
363 1220
363 1258
348 1258
1 1 2 0 0 0 0 146 148 0 0 3
168 1242
278 1242
278 1249
3 0 85 0 0 0 0 148 0 0 305 2
272 1267
262 1267
0 2 85 0 0 28800 0 0 148 158 0 12
2200 1470
2181 1470
2181 1659
1657 1659
1657 2247
1880 2247
1880 2601
50 2601
50 1307
262 1307
262 1258
272 1258
0 4 90 0 0 0 0 0 148 334 0 3
102 1001
102 1276
278 1276
0 5 65 0 0 0 0 0 148 335 0 5
776 1083
776 1160
200 1160
200 1285
278 1285
0 6 64 0 0 0 0 0 148 336 0 5
803 1074
803 1180
214 1180
214 1294
278 1294
0 7 45 0 0 8320 0 0 148 337 0 5
829 1064
829 1189
228 1189
228 1303
278 1303
0 8 63 0 0 8320 0 0 148 338 0 5
855 1056
855 1210
247 1210
247 1312
278 1312
1 0 63 0 0 0 0 149 0 0 338 2
666 1041
855 1041
1 0 45 0 0 0 0 150 0 0 337 2
646 1031
829 1031
1 0 64 0 0 0 0 151 0 0 336 2
625 1023
803 1023
1 0 65 0 0 0 0 152 0 0 335 2
597 1015
776 1015
14 1 63 0 0 0 0 158 149 0 0 3
547 1040
547 1041
666 1041
13 1 45 0 0 0 0 158 150 0 0 2
547 1031
646 1031
12 1 64 0 0 0 0 158 151 0 0 3
547 1022
547 1023
625 1023
11 1 65 0 0 0 0 158 152 0 0 3
547 1013
547 1015
597 1015
1 0 2 0 0 0 0 158 0 0 320 3
483 977
483 898
387 898
1 0 2 0 0 0 0 159 0 0 321 4
289 977
289 898
388 898
388 977
9 0 2 0 0 0 0 159 0 0 322 3
359 977
388 977
388 986
10 1 2 0 0 0 0 159 153 0 0 3
359 986
388 986
388 992
9 0 86 0 0 4096 0 158 0 0 324 4
553 977
576 977
576 998
553 998
10 0 86 0 0 24704 0 158 0 0 159 13
553 986
553 1169
77 1169
77 1117
44 1117
44 2606
1886 2606
1886 2239
1670 2239
1670 1646
2100 1646
2100 1469
2119 1469
2 0 87 0 0 0 0 158 0 0 326 2
477 986
468 986
0 3 87 0 0 8192 0 0 158 328 0 5
263 987
263 948
468 948
468 995
477 995
3 0 87 0 0 0 0 159 0 0 328 2
283 995
263 995
0 2 87 0 0 28800 0 0 159 160 0 12
2047 1470
2016 1470
2016 1636
1683 1636
1683 2229
1893 2229
1893 2610
40 2610
40 1058
263 1058
263 986
283 986
11 1 40 0 0 0 0 159 157 0 0 6
353 1013
368 1013
368 1063
276 1063
276 1145
302 1145
12 1 43 0 0 0 0 159 156 0 0 5
353 1022
353 1077
323 1077
323 1144
337 1144
13 1 41 0 0 0 0 159 155 0 0 4
353 1031
360 1031
360 1142
374 1142
14 1 42 0 0 0 0 159 154 0 0 4
353 1040
403 1040
403 1147
419 1147
0 4 90 0 0 0 0 0 158 334 0 5
235 1001
235 917
453 917
453 1004
483 1004
0 4 90 0 0 0 0 0 159 387 0 6
257 393
102 393
102 1001
235 1001
235 1004
289 1004
0 5 65 0 0 0 0 0 158 354 0 5
776 833
776 1084
454 1084
454 1013
483 1013
0 6 64 0 0 0 0 0 158 353 0 5
803 842
803 1075
463 1075
463 1022
483 1022
0 7 45 0 0 0 0 0 158 352 0 5
829 851
829 1065
474 1065
474 1031
483 1031
0 8 63 0 0 0 0 0 158 351 0 4
855 860
855 1057
483 1057
483 1040
0 8 123 0 0 8192 0 0 159 355 0 5
743 823
743 943
173 943
173 1040
289 1040
0 7 124 0 0 8192 0 0 159 356 0 5
719 815
719 935
187 935
187 1031
289 1031
0 6 125 0 0 8192 0 0 159 357 0 5
694 805
694 925
198 925
198 1022
289 1022
0 5 126 0 0 8192 0 0 159 358 0 5
667 795
667 908
213 908
213 1013
289 1013
1 0 63 0 0 0 0 161 0 0 351 2
850 862
850 860
1 0 45 0 0 0 0 162 0 0 352 2
822 851
822 851
1 0 64 0 0 0 0 163 0 0 353 2
790 844
790 842
1 0 65 0 0 0 0 164 0 0 354 2
763 835
763 833
1 0 123 0 0 0 0 165 0 0 355 2
733 825
733 824
1 0 124 0 0 0 0 166 0 0 356 2
712 817
712 815
1 0 125 0 0 0 0 167 0 0 357 2
681 806
681 806
1 0 126 0 0 0 0 168 0 0 358 2
639 797
639 797
0 18 63 0 0 0 0 0 170 391 0 3
855 463
855 860
519 860
0 17 45 0 0 0 0 0 170 390 0 3
829 482
829 851
519 851
0 16 64 0 0 0 0 0 170 389 0 3
803 503
803 842
519 842
0 15 65 0 0 0 0 0 170 388 0 3
776 525
776 833
519 833
0 14 123 0 0 4224 0 0 170 0 0 3
743 69
743 824
519 824
0 13 124 0 0 4224 0 0 170 0 0 3
719 70
719 815
519 815
0 12 125 0 0 4224 0 0 170 0 0 5
695 70
695 805
694 805
694 806
519 806
0 11 126 0 0 4224 0 0 170 0 0 5
668 72
668 795
667 795
667 797
519 797
1 0 127 0 0 4096 0 173 0 0 360 2
556 586
556 605
12 9 127 0 0 12416 0 176 170 0 0 6
520 605
557 605
557 708
407 708
407 851
455 851
20 1 128 0 0 4224 0 170 160 0 0 3
525 788
597 788
597 767
0 19 3 0 0 28800 0 0 170 161 0 13
1974 1469
1964 1469
1964 1626
1693 1626
1693 2221
1897 2221
1897 2616
36 2616
36 763
338 763
338 738
525 738
525 779
1 0 129 0 0 4096 0 170 0 0 368 2
455 779
443 779
2 0 129 0 0 0 0 170 0 0 368 2
455 788
443 788
3 0 129 0 0 0 0 170 0 0 368 2
455 797
443 797
4 0 129 0 0 0 0 170 0 0 368 2
455 806
443 806
5 0 129 0 0 0 0 170 0 0 368 2
455 815
443 815
0 6 129 0 0 4224 0 0 170 0 0 4
373 773
443 773
443 824
455 824
0 7 130 0 0 8320 0 0 170 372 0 5
604 641
604 730
436 730
436 833
455 833
0 8 131 0 0 8320 0 0 170 373 0 5
583 623
583 718
419 718
419 842
455 842
1 10 132 0 0 12416 0 174 170 0 0 5
532 588
532 698
394 698
394 860
455 860
14 1 130 0 0 0 0 176 171 0 0 3
520 641
604 641
604 584
13 1 131 0 0 0 0 176 172 0 0 3
520 623
583 623
583 582
11 1 132 0 0 0 0 176 174 0 0 3
520 587
520 588
532 588
1 10 2 0 0 0 0 175 176 0 0 3
430 678
430 650
450 650
1 8 133 0 0 12416 0 19 176 0 0 4
279 710
365 710
365 632
456 632
1 6 134 0 0 12416 0 20 176 0 0 4
282 656
340 656
340 614
456 614
1 4 135 0 0 4224 0 21 176 0 0 4
282 607
374 607
374 596
456 596
1 2 136 0 0 12416 0 22 176 0 0 4
284 557
328 557
328 578
456 578
1 1 137 0 0 12416 0 23 176 0 0 6
227 536
237 536
237 506
383 506
383 569
456 569
11 9 138 0 0 12416 0 177 176 0 0 6
527 406
588 406
588 470
394 470
394 641
456 641
12 7 139 0 0 12416 0 177 176 0 0 6
527 415
573 415
573 493
413 493
413 623
456 623
13 5 140 0 0 12416 0 177 176 0 0 6
527 424
553 424
553 514
433 514
433 605
456 605
14 3 141 0 0 8320 0 177 176 0 0 6
527 433
535 433
535 537
442 537
442 587
456 587
3 0 88 0 0 4096 0 177 0 0 386 4
457 388
403 388
403 384
388 384
0 2 88 0 0 32896 0 0 177 162 0 12
1902 1470
1889 1470
1889 1611
1704 1611
1704 2210
1904 2210
1904 2621
27 2621
27 463
388 463
388 379
457 379
4 0 90 0 0 0 0 177 0 0 412 3
463 397
257 397
257 63
0 5 65 0 0 0 0 0 177 395 0 5
776 223
776 526
403 526
403 406
463 406
0 6 64 0 0 0 0 0 177 396 0 5
803 243
803 503
423 503
423 415
463 415
0 7 45 0 0 0 0 0 177 397 0 5
829 266
829 483
443 483
443 424
463 424
0 8 63 0 0 0 0 0 177 398 0 4
855 293
855 463
463 463
463 433
10 0 2 0 0 0 0 177 0 0 393 3
533 379
543 379
543 366
9 0 2 0 0 0 0 177 0 0 394 5
533 370
543 370
543 323
442 323
442 366
1 1 2 0 0 0 0 178 177 0 0 7
323 177
323 165
296 165
296 366
442 366
442 370
463 370
0 5 65 0 0 0 0 0 180 399 0 5
776 88
776 223
370 223
370 115
394 115
0 6 64 0 0 0 0 0 180 400 0 5
803 106
803 243
380 243
380 124
394 124
0 7 45 0 0 0 0 0 180 401 0 5
829 124
829 267
388 267
388 133
394 133
0 8 63 0 0 0 0 0 180 402 0 4
855 142
855 293
394 293
394 142
9 0 65 0 0 0 0 179 0 0 0 5
620 88
776 88
776 88
775 88
775 67
10 0 64 0 0 0 0 179 0 0 0 5
620 106
803 106
803 106
802 106
802 67
11 0 45 0 0 0 0 179 0 0 0 5
620 124
829 124
829 124
828 124
828 68
12 0 63 0 0 0 0 179 0 0 0 5
620 142
855 142
855 142
853 142
853 67
0 7 27 0 0 0 0 0 179 404 0 3
542 115
542 133
556 133
0 5 27 0 0 0 0 0 179 405 0 3
538 97
538 115
556 115
0 3 27 0 0 0 0 0 179 406 0 3
538 79
538 97
556 97
1 0 27 0 0 32896 0 179 0 0 0 16
556 79
538 79
538 20
34 20
34 370
77 370
77 407
13 407
13 2637
1920 2637
1920 2191
1736 2191
1736 1577
1791 1577
1791 1470
1806 1470
3 0 83 0 0 16512 0 180 0 0 154 12
388 97
77 97
77 305
20 305
20 2631
1913 2631
1913 2200
1719 2200
1719 1593
2396 1593
2396 1459
2421 1459
11 2 82 0 0 12416 0 180 179 0 0 4
458 115
485 115
485 88
556 88
12 4 81 0 0 12416 0 180 179 0 0 4
458 124
502 124
502 106
556 106
13 6 80 0 0 4224 0 180 179 0 0 4
458 133
512 133
512 124
556 124
14 8 79 0 0 4224 0 180 179 0 0 2
458 142
556 142
3 1 90 0 0 0 0 181 180 0 0 3
200 63
394 63
394 79
0 2 142 0 0 4224 0 0 181 0 0 3
145 76
145 72
146 72
1 1 143 0 0 4224 0 181 24 0 0 4
152 63
118 63
118 71
105 71
45
-24 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
946 2366 1053 2407
957 2374 1041 2401
6 output
-24 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
929 1329 968 1370
941 1338 955 1365
1 z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1043 1430 1094 1454
1054 1438 1082 1454
4 cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2565 1505 2584 1521
2565 1505 2584 1521
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2496 1509 2515 1525
2496 1509 2515 1525
2 EB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2414 1513 2433 1529
2414 1513 2433 1529
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2336 1513 2355 1529
2336 1513 2355 1529
2 Lo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2261 1524 2280 1540
2261 1524 2280 1540
2 EA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2191 1512 2210 1528
2191 1512 2210 1528
2 LA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2112 1516 2131 1532
2112 1516 2131 1532
2 Ei
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
2038 1516 2057 1532
2038 1516 2057 1532
2 Li
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1965 1514 1984 1530
1965 1514 1984 1530
2 CE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1892 1515 1911 1531
1892 1515 1911 1531
2 LM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1813 1518 1832 1534
1813 1518 1832 1534
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1732 1519 1751 1535
1732 1519 1751 1535
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1704 548 1723 564
1704 548 1723 564
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1704 490 1723 506
1704 490 1723 506
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1696 421 1715 437
1696 421 1715 437
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1677 362 1696 378
1677 362 1696 378
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1318 78 1357 102
1330 87 1344 103
2 I4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1262 80 1299 104
1273 88 1287 104
2 I5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1213 75 1250 99
1224 84 1238 100
2 I6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1163 76 1200 100
1174 85 1188 101
2 I7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
535 2220 612 2242
545 2227 601 2243
7 O/P REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
290 2178 349 2199
299 2184 339 2199
5 C REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
553 2112 596 2133
562 2118 586 2133
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
478 1701 537 1722
487 1707 527 1722
5 B REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
534 1547 575 1568
542 1553 566 1568
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
148 1385 191 1406
157 1392 181 1407
3 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
147 1413 196 1434
155 1420 187 1435
4 mode
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
212 1476 245 1497
220 1482 236 1497
2 s0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
212 1451 247 1472
221 1457 237 1472
2 s1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
212 1425 247 1446
221 1431 237 1446
2 s2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
212 1399 247 1420
221 1406 237 1421
2 s3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
380 1221 485 1242
388 1228 476 1243
11 ACCUMULATOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
726 -2 785 19
735 4 775 19
5 W BUS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
60 21 165 42
68 28 156 43
11 CLOCK PULSE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
389 1005 422 1026
397 1011 413 1026
2 IR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
527 754 570 775
536 761 560 776
3 RAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
469 662 512 683
478 669 502 684
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
593 373 636 394
602 379 626 394
3 MAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
189 610 248 631
198 617 238 632
5 INPUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
489 141 524 162
498 148 514 163
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1004 7 1034 31
1015 16 1022 32
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1681 177 1786 198
1689 184 1777 199
11 CLOCK PULSE
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
