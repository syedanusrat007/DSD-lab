CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
52
13 Logic Switch~
5 276 573 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
3 V36
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5433 0 0
2
42919 0
0
13 Logic Switch~
5 254 565 0 1 11
0 7
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V35
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3679 0 0
2
42919 0
0
13 Logic Switch~
5 226 556 0 1 11
0 8
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V34
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9342 0 0
2
42919 0
0
13 Logic Switch~
5 203 549 0 1 11
0 9
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V33
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3623 0 0
2
42919 0
0
13 Logic Switch~
5 183 538 0 1 11
0 10
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V32
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3722 0 0
2
42919 0
0
13 Logic Switch~
5 159 529 0 1 11
0 11
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V31
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8993 0 0
2
42919 0
0
13 Logic Switch~
5 137 520 0 1 11
0 12
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V30
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3723 0 0
2
42919 0
0
13 Logic Switch~
5 115 511 0 1 11
0 13
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V29
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6244 0 0
2
42919 0
0
13 Logic Switch~
5 277 449 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
3 V28
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6421 0 0
2
42919 0
0
13 Logic Switch~
5 248 440 0 1 11
0 15
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V27
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7743 0 0
2
42919 0
0
13 Logic Switch~
5 224 431 0 1 11
0 16
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9840 0 0
2
42919 0
0
13 Logic Switch~
5 203 421 0 1 11
0 17
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V25
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6910 0 0
2
42919 0
0
13 Logic Switch~
5 183 414 0 1 11
0 18
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V24
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
449 0 0
2
42919 0
0
13 Logic Switch~
5 162 404 0 1 11
0 19
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V23
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8761 0 0
2
42919 0
0
13 Logic Switch~
5 134 395 0 1 11
0 20
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6748 0 0
2
42919 0
0
13 Logic Switch~
5 115 386 0 1 11
0 21
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7393 0 0
2
42919 0
0
13 Logic Switch~
5 274 319 0 1 11
0 22
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7699 0 0
2
42919 0
0
13 Logic Switch~
5 247 310 0 1 11
0 23
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6638 0 0
2
42919 0
0
13 Logic Switch~
5 221 301 0 1 11
0 24
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4595 0 0
2
42919 0
0
13 Logic Switch~
5 201 292 0 1 11
0 25
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9395 0 0
2
42919 0
0
13 Logic Switch~
5 177 283 0 1 11
0 26
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3303 0 0
2
42919 0
0
13 Logic Switch~
5 154 275 0 1 11
0 27
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4498 0 0
2
42919 0
0
13 Logic Switch~
5 136 264 0 1 11
0 28
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9728 0 0
2
42919 0
0
13 Logic Switch~
5 116 256 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3789 0 0
2
42919 0
0
13 Logic Switch~
5 90 112 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3978 0 0
2
42919 0
0
13 Logic Switch~
5 275 176 0 1 11
0 31
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3494 0 0
2
42919 0
0
13 Logic Switch~
5 246 166 0 1 11
0 32
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3507 0 0
2
42919 0
0
13 Logic Switch~
5 221 158 0 1 11
0 33
0
0 0 21360 692
2 0V
-7 -16 7 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5151 0 0
2
42919 0
0
13 Logic Switch~
5 203 147 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3701 0 0
2
42919 0
0
13 Logic Switch~
5 173 139 0 1 11
0 35
0
0 0 21360 692
2 0V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8585 0 0
2
42919 0
0
13 Logic Switch~
5 147 130 0 1 11
0 36
0
0 0 21360 692
2 0V
-7 -16 7 -8
2 V7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8809 0 0
2
42919 0
0
13 Logic Switch~
5 120 121 0 1 11
0 37
0
0 0 21360 692
2 0V
-7 -16 7 -8
2 V6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5993 0 0
2
42919 0
0
13 Logic Switch~
5 776 132 0 1 11
0 2
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V4
-1 -24 13 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8654 0 0
2
42919 0
0
13 Logic Switch~
5 814 89 0 1 11
0 3
0
0 0 21360 512
2 0V
0 -16 14 -8
2 V3
4 -22 18 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7223 0 0
2
42919 0
0
13 Logic Switch~
5 797 54 0 1 11
0 4
0
0 0 21360 512
2 0V
24 -17 38 -9
2 V2
-1 -24 13 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3641 0 0
2
42919 0
0
13 Logic Switch~
5 880 33 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V1
29 -24 43 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3104 0 0
2
42919 0
0
14 Logic Display~
6 896 588 0 1 2
10 44
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3296 0 0
2
42919 0
0
14 Logic Display~
6 897 561 0 1 2
10 45
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8534 0 0
2
42919 0
0
14 Logic Display~
6 900 472 0 1 2
10 38
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
949 0 0
2
42919 0
0
14 Logic Display~
6 897 436 0 1 2
10 39
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3371 0 0
2
42919 0
0
14 Logic Display~
6 902 334 0 1 2
10 40
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7311 0 0
2
42919 0
0
14 Logic Display~
6 901 306 0 1 2
10 41
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
42919 0
0
14 Logic Display~
6 909 185 0 1 2
10 42
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3526 0 0
2
42919 0
0
14 Logic Display~
6 902 162 0 1 2
10 43
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4129 0 0
2
42919 0
0
9 Inverter~
13 693 132 0 2 22
0 2 46
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U5D
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6278 0 0
2
42919 0
0
9 Inverter~
13 748 89 0 2 22
0 3 47
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U5C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3482 0 0
2
42919 0
0
9 Inverter~
13 725 54 0 2 22
0 4 48
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U5B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8323 0 0
2
42919 0
0
9 Inverter~
13 802 34 0 2 22
0 5 49
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U5A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3984 0 0
2
42919 0
0
7 74LS151
20 347 538 0 14 29
0 13 12 11 10 9 8 7 6 49
48 47 46 45 44
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
7622 0 0
2
42919 0
0
7 74LS151
20 349 413 0 14 29
0 21 50 19 18 17 16 15 14 49
48 47 46 39 38
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
816 0 0
2
42919 0
0
7 74LS151
20 350 283 0 14 29
0 29 28 27 26 25 24 23 22 49
48 47 46 41 40
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
4656 0 0
2
42919 0
0
7 74LS151
20 352 139 0 14 29
0 30 37 36 35 34 33 32 31 49
48 47 46 43 42
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
6356 0 0
2
42919 0
0
109
1 0 2 0 0 4096 0 33 0 0 2 2
764 132
717 132
1 1 2 0 0 4224 0 45 33 0 0 2
714 132
764 132
1 1 2 0 0 0 0 33 45 0 0 2
764 132
714 132
1 0 3 0 0 4096 0 34 0 0 83 2
802 89
772 89
0 1 4 0 0 4096 0 0 35 6 0 2
751 54
785 54
1 0 4 0 0 0 0 35 0 0 0 4
785 54
751 54
751 54
755 54
0 1 5 0 0 4096 0 0 36 73 0 2
826 33
868 33
1 0 6 0 0 4096 0 1 0 0 41 2
288 573
288 574
1 0 7 0 0 0 0 2 0 0 44 2
266 565
266 565
1 0 8 0 0 0 0 3 0 0 47 2
238 556
238 556
1 0 9 0 0 4096 0 4 0 0 50 2
215 549
215 547
1 0 10 0 0 0 0 5 0 0 53 2
195 538
195 538
1 0 11 0 0 0 0 6 0 0 56 2
171 529
171 529
1 0 12 0 0 0 0 7 0 0 59 2
149 520
149 520
1 0 13 0 0 0 0 8 0 0 62 2
127 511
127 511
1 0 14 0 0 0 0 9 0 0 42 2
289 449
289 449
1 0 15 0 0 0 0 10 0 0 45 2
260 440
260 440
1 0 16 0 0 0 0 11 0 0 48 2
236 431
236 431
1 0 17 0 0 4096 0 12 0 0 51 2
215 421
215 422
1 0 18 0 0 4096 0 13 0 0 54 2
195 414
195 413
1 0 19 0 0 0 0 14 0 0 57 2
174 404
174 404
1 0 20 0 0 0 0 15 0 0 60 2
146 395
146 395
1 0 21 0 0 0 0 16 0 0 63 2
127 386
127 386
1 0 22 0 0 0 0 17 0 0 43 2
286 319
286 319
1 0 23 0 0 0 0 18 0 0 46 2
259 310
259 310
1 0 24 0 0 0 0 19 0 0 49 2
233 301
233 301
1 0 25 0 0 0 0 20 0 0 52 2
213 292
213 292
1 0 26 0 0 0 0 21 0 0 55 2
189 283
189 283
1 0 27 0 0 4096 0 22 0 0 58 2
166 275
166 274
1 0 28 0 0 4096 0 23 0 0 61 2
148 264
148 265
1 0 29 0 0 0 0 24 0 0 64 2
128 256
128 256
1 0 30 0 0 0 0 25 0 0 33 2
102 112
102 112
0 0 30 0 0 4096 0 0 0 0 72 2
83 112
137 112
1 0 31 0 0 4096 0 26 0 0 65 2
287 176
287 175
1 0 32 0 0 0 0 27 0 0 66 2
258 166
258 166
1 0 33 0 0 4096 0 28 0 0 67 2
233 158
233 157
1 0 34 0 0 4096 0 29 0 0 68 2
215 147
215 148
1 0 35 0 0 0 0 30 0 0 69 2
185 139
185 139
1 0 36 0 0 0 0 31 0 0 70 2
159 130
159 130
1 0 37 0 0 0 0 32 0 0 71 2
132 121
132 121
8 0 6 0 0 4224 0 49 0 0 0 2
315 574
267 574
8 0 14 0 0 4224 0 50 0 0 0 2
317 449
267 449
8 0 22 0 0 4224 0 51 0 0 0 2
318 319
266 319
7 0 7 0 0 4224 0 49 0 0 0 2
315 565
242 565
7 0 15 0 0 4224 0 50 0 0 0 2
317 440
241 440
7 0 23 0 0 4224 0 51 0 0 0 2
318 310
241 310
6 0 8 0 0 4224 0 49 0 0 0 2
315 556
213 556
6 0 16 0 0 4224 0 50 0 0 0 2
317 431
212 431
6 0 24 0 0 4224 0 51 0 0 0 2
318 301
211 301
5 0 9 0 0 4224 0 49 0 0 0 2
315 547
194 547
5 0 17 0 0 4224 0 50 0 0 0 2
317 422
192 422
5 0 25 0 0 4224 0 51 0 0 0 2
318 292
192 292
4 0 10 0 0 4224 0 49 0 0 0 2
315 538
170 538
4 0 18 0 0 4224 0 50 0 0 0 2
317 413
170 413
4 0 26 0 0 4224 0 51 0 0 0 2
318 283
167 283
3 0 11 0 0 4224 0 49 0 0 0 2
315 529
146 529
3 0 19 0 0 4224 0 50 0 0 0 2
317 404
146 404
3 0 27 0 0 4224 0 51 0 0 0 2
318 274
145 274
2 0 12 0 0 4224 0 49 0 0 0 2
315 520
124 520
0 0 20 0 0 4224 0 0 0 0 0 2
323 395
124 395
2 0 28 0 0 4224 0 51 0 0 0 2
318 265
125 265
1 0 13 0 0 4224 0 49 0 0 0 2
315 511
113 511
1 0 21 0 0 4224 0 50 0 0 0 2
317 386
112 386
1 0 29 0 0 4224 0 51 0 0 0 2
318 256
112 256
8 0 31 0 0 4224 0 52 0 0 0 2
320 175
266 175
7 0 32 0 0 4224 0 52 0 0 0 2
320 166
239 166
6 0 33 0 0 4224 0 52 0 0 0 2
320 157
210 157
5 0 34 0 0 4224 0 52 0 0 0 2
320 148
188 148
4 0 35 0 0 4224 0 52 0 0 0 2
320 139
165 139
3 0 36 0 0 4224 0 52 0 0 0 2
320 130
144 130
2 0 37 0 0 4224 0 52 0 0 0 2
320 121
124 121
1 0 30 0 0 4224 0 52 0 0 0 2
320 112
112 112
1 0 5 0 0 0 0 36 0 0 0 4
868 33
826 33
826 34
830 34
1 0 38 0 0 4096 0 39 0 0 105 2
884 476
863 476
1 0 39 0 0 4096 0 40 0 0 106 2
881 440
872 440
1 0 40 0 0 8192 0 41 0 0 103 3
886 338
886 337
861 337
1 0 41 0 0 4096 0 42 0 0 104 2
885 310
869 310
1 0 42 0 0 4096 0 43 0 0 101 2
893 189
875 189
1 0 43 0 0 4096 0 44 0 0 102 2
886 166
872 166
1 0 44 0 0 0 0 37 0 0 107 2
880 592
880 592
1 0 45 0 0 0 0 38 0 0 108 2
881 565
881 565
1 1 2 0 0 0 0 33 45 0 0 2
764 132
714 132
1 1 3 0 0 4224 0 34 46 0 0 2
802 89
769 89
1 1 4 0 0 4224 0 35 47 0 0 2
785 54
746 54
1 1 5 0 0 4224 0 36 48 0 0 4
868 33
822 33
822 34
823 34
12 0 46 0 0 4096 0 51 0 0 88 2
382 283
578 283
12 0 46 0 0 4096 0 50 0 0 88 2
381 413
578 413
0 12 46 0 0 4224 0 0 49 109 0 3
578 132
578 538
379 538
11 0 47 0 0 4096 0 51 0 0 91 2
382 274
534 274
11 0 47 0 0 4096 0 50 0 0 91 2
381 404
534 404
0 11 47 0 0 4224 0 0 49 100 0 3
534 89
534 529
379 529
10 0 48 0 0 4096 0 51 0 0 94 2
382 265
489 265
10 0 48 0 0 4096 0 50 0 0 94 2
381 395
489 395
0 10 48 0 0 4224 0 0 49 99 0 3
489 53
489 520
379 520
9 0 49 0 0 4096 0 51 0 0 97 2
388 256
445 256
9 0 49 0 0 4096 0 50 0 0 97 2
387 386
445 386
0 9 49 0 0 4224 0 0 49 98 0 3
445 34
445 511
385 511
9 2 49 0 0 128 0 52 48 0 0 3
390 112
390 34
787 34
10 2 48 0 0 128 0 52 47 0 0 4
384 121
384 53
710 53
710 54
11 2 47 0 0 128 0 52 46 0 0 3
384 130
384 89
733 89
14 1 42 0 0 8320 0 52 43 0 0 3
390 175
390 189
893 189
13 1 43 0 0 4224 0 52 44 0 0 2
384 166
886 166
14 1 40 0 0 8320 0 51 41 0 0 4
388 319
388 337
886 337
886 338
13 1 41 0 0 4224 0 51 42 0 0 2
382 310
885 310
14 1 38 0 0 8320 0 50 39 0 0 3
387 449
387 476
884 476
13 1 39 0 0 4224 0 50 40 0 0 2
381 440
881 440
14 0 44 0 0 8320 0 49 0 0 0 3
385 574
385 592
886 592
13 0 45 0 0 4224 0 49 0 0 0 2
379 565
885 565
12 2 46 0 0 128 0 52 45 0 0 3
384 139
384 132
678 132
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
