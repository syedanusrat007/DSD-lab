CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
290 1260 15 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
132
13 Logic Switch~
5 206 441 0 10 11
0 85 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
42999.8 0
0
13 Logic Switch~
5 321 1462 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V31
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89816e-315 0
0
13 Logic Switch~
5 380 501 0 10 11
0 86 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V20
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89816e-315 5.26354e-315
0
13 Logic Switch~
5 348 500 0 1 11
0 87
0
0 0 21360 90
2 0V
11 0 25 8
3 V22
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89816e-315 5.30499e-315
0
13 Logic Switch~
5 317 500 0 1 11
0 88
0
0 0 21360 90
2 0V
11 0 25 8
3 V23
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89816e-315 5.32571e-315
0
13 Logic Switch~
5 284 498 0 1 11
0 89
0
0 0 21360 90
2 0V
11 0 25 8
3 V24
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89816e-315 5.34643e-315
0
13 Logic Switch~
5 1536 965 0 1 11
0 110
0
0 0 21360 90
2 0V
11 0 25 8
3 V12
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89816e-315 5.3568e-315
0
13 Logic Switch~
5 1569 967 0 1 11
0 109
0
0 0 21360 90
2 0V
11 0 25 8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.89816e-315 5.36716e-315
0
13 Logic Switch~
5 1600 967 0 1 11
0 108
0
0 0 21360 90
2 0V
11 0 25 8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.89816e-315 5.37752e-315
0
13 Logic Switch~
5 1632 968 0 10 11
0 107 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.89816e-315 5.38788e-315
0
13 Logic Switch~
5 1385 966 0 10 11
0 98 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.89816e-315 5.39306e-315
0
13 Logic Switch~
5 1353 965 0 1 11
0 97
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.89816e-315 5.39824e-315
0
13 Logic Switch~
5 1322 965 0 1 11
0 96
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
5.89816e-315 5.40342e-315
0
13 Logic Switch~
5 1289 963 0 1 11
0 95
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.89816e-315 5.4086e-315
0
14 Logic Display~
6 1621 744 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L53
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
43000.7 0
0
14 Logic Display~
6 1577 1014 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L52
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
43000.7 0
0
14 Logic Display~
6 416 1057 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L51
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
43000.7 0
0
9 2-In AND~
219 939 1770 0 3 22
0 39 7 6
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U30D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
9323 0 0
2
5.89816e-315 0
0
5 4025~
219 851 1718 0 4 22
0 24 8 10 25
0
0 0 624 270
4 4025
-14 -24 14 -16
4 U32A
32 -10 60 -2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 15 0
1 U
317 0 0
2
42999.8 1
0
8 2-In OR~
219 574 1703 0 3 22
0 10 8 9
0
0 0 624 180
5 74F32
-18 -24 17 -16
4 U26B
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3108 0 0
2
42999.8 2
0
9 2-In AND~
219 630 1694 0 3 22
0 11 12 8
0
0 0 624 180
5 74F08
-18 -24 17 -16
4 U30C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
4299 0 0
2
42999.8 3
0
14 Logic Display~
6 1088 945 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L50
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89816e-315 5.41378e-315
0
14 Logic Display~
6 1114 948 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L49
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89816e-315 5.41896e-315
0
14 Logic Display~
6 1139 947 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L37
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89816e-315 5.42414e-315
0
14 Logic Display~
6 1163 947 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L36
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89816e-315 5.42933e-315
0
14 Logic Display~
6 382 1871 0 1 2
10 17
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L48
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89816e-315 5.43192e-315
0
14 Logic Display~
6 462 1879 0 1 2
10 17
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L47
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89816e-315 5.43451e-315
0
14 Logic Display~
6 488 1878 0 1 2
10 9
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L46
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89816e-315 5.4371e-315
0
14 Logic Display~
6 1431 1911 0 1 2
10 23
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L45
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89816e-315 5.43969e-315
0
14 Logic Display~
6 1399 1908 0 1 2
10 22
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L44
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89816e-315 5.44228e-315
0
14 Logic Display~
6 1367 1915 0 1 2
10 21
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L43
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89816e-315 5.44487e-315
0
14 Logic Display~
6 1341 1918 0 1 2
10 20
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L42
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.89816e-315 5.44746e-315
0
14 Logic Display~
6 1300 1920 0 1 2
10 19
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L41
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.89816e-315 5.45005e-315
0
14 Logic Display~
6 1259 1927 0 1 2
10 18
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89816e-315 5.45264e-315
0
14 Logic Display~
6 920 1905 0 1 2
10 6
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L39
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.89816e-315 5.45523e-315
0
14 Logic Display~
6 633 1886 0 1 2
10 24
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L38
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.89816e-315 5.45782e-315
0
14 Logic Display~
6 822 1872 0 1 2
10 25
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L35
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89816e-315 5.46041e-315
0
14 Logic Display~
6 667 1844 0 1 2
10 7
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L34
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89816e-315 5.463e-315
0
9 2-In AND~
219 337 1200 0 3 22
0 27 13 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U30B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
9281 0 0
2
42999.8 4
0
9 2-In XOR~
219 386 1369 0 3 22
0 2 10 28
0
0 0 624 90
6 74LS86
-21 -24 21 -16
4 U31A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
8464 0 0
2
5.89816e-315 5.46559e-315
0
7 Ground~
168 380 1392 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
5.89816e-315 5.46818e-315
0
7 Ground~
168 571 1263 0 1 3
0 2
0
0 0 53360 180
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
5.89816e-315 5.47077e-315
0
9 Inverter~
13 1776 762 0 2 22
0 22 3
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U29C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
4139 0 0
2
42999.8 5
0
9 2-In NOR~
219 939 1714 0 3 22
0 52 17 39
0
0 0 624 270
4 7428
-14 -24 14 -16
4 U28C
32 -10 60 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
6435 0 0
2
42999.8 6
0
9 Inverter~
13 1699 1031 0 2 22
0 18 4
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U29B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
5283 0 0
2
5.89816e-315 5.47207e-315
0
9 2-In NOR~
219 990 1818 0 3 22
0 59 52 19
0
0 0 624 270
4 7428
-14 -24 14 -16
4 U28B
32 -10 60 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
6874 0 0
2
5.89816e-315 5.47336e-315
0
9 Inverter~
13 320 1059 0 2 22
0 17 5
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U29A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
5305 0 0
2
5.89816e-315 5.47466e-315
0
5 4011~
219 740 1752 0 3 22
0 54 12 7
0
0 0 624 180
4 4011
-7 -24 21 -16
4 U27A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 10 0
1 U
34 0 0
2
5.89816e-315 5.47595e-315
0
9 Inverter~
13 1854 587 0 2 22
0 23 76
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U19F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
969 0 0
2
42999.8 7
0
9 Inverter~
13 1852 545 0 2 22
0 22 75
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U19E
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
8402 0 0
2
42999.8 8
0
9 2-In AND~
219 1095 1787 0 3 22
0 54 53 21
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3751 0 0
2
42999.8 9
0
9 2-In AND~
219 1185 1744 0 3 22
0 55 54 20
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
4292 0 0
2
42999.8 10
0
9 2-In AND~
219 1127 1689 0 3 22
0 54 56 18
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6118 0 0
2
42999.8 11
0
8 2-In OR~
219 1039 1696 0 3 22
0 55 53 57
0
0 0 624 270
5 74F32
-18 -24 17 -16
4 U26A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
34 0 0
2
42999.8 12
0
8 3-In OR~
219 1029 1640 0 4 22
0 58 22 23 53
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U25A
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
6357 0 0
2
42999.8 13
0
9 2-In AND~
219 1026 1765 0 3 22
0 57 54 59
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
319 0 0
2
42999.8 14
0
9 2-In AND~
219 957 1666 0 3 22
0 60 11 52
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3976 0 0
2
42999.8 15
0
9 2-In AND~
219 877 1662 0 3 22
0 54 60 24
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7634 0 0
2
42999.8 16
0
8 2-In OR~
219 770 1702 0 3 22
0 62 61 12
0
0 0 624 270
5 74F32
-18 -24 17 -16
4 U23A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
523 0 0
2
42999.8 17
0
9 2-In AND~
219 784 1661 0 3 22
0 29 63 62
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6748 0 0
2
42999.8 18
0
2 +V
167 675 1372 0 1 3
0 64
0
0 0 54256 180
3 10V
6 -2 27 6
3 V32
6 -12 27 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6901 0 0
2
42999.8 19
0
9 3-In NOR~
219 711 1261 0 4 22
0 10 17 54 65
0
0 0 624 180
5 74F27
-18 -24 17 -16
4 U21A
-11 -2 17 6
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
842 0 0
2
42999.8 20
0
14 Logic Display~
6 1552 1300 0 1 2
10 54
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L33
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
42999.8 21
0
14 Logic Display~
6 1552 1325 0 1 2
10 17
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L32
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
42999.8 22
0
14 Logic Display~
6 1552 1351 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L31
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
42999.8 23
0
14 Logic Display~
6 1552 1274 0 1 2
10 11
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L30
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
42999.8 24
0
7 74LS164
127 716 1324 0 12 25
0 65 65 26 64 111 112 113 114 11
54 17 10
0
0 0 4848 0
6 74F164
-21 -51 21 -43
3 U20
-14 4 7 12
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
6986 0 0
2
42999.8 25
0
14 Logic Display~
6 1550 1405 0 1 2
10 60
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L21
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
5.89816e-315 5.47725e-315
0
14 Logic Display~
6 1550 1482 0 1 2
10 58
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L23
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
5.89816e-315 5.47854e-315
0
14 Logic Display~
6 1550 1456 0 1 2
10 22
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L24
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.89816e-315 5.47984e-315
0
14 Logic Display~
6 1549 1558 0 1 2
10 61
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L25
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89816e-315 5.48113e-315
0
14 Logic Display~
6 1550 1584 0 1 2
10 63
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L26
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
5.89816e-315 5.48243e-315
0
14 Logic Display~
6 1549 1533 0 1 2
10 56
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L27
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9466 0 0
2
5.89816e-315 5.48372e-315
0
14 Logic Display~
6 1549 1507 0 1 2
10 55
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L28
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3266 0 0
2
5.89816e-315 5.48502e-315
0
14 Logic Display~
6 1550 1608 0 1 2
10 66
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L29
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
5.89816e-315 5.48631e-315
0
14 Logic Display~
6 1550 1431 0 1 2
10 23
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3723 0 0
2
5.89816e-315 5.48761e-315
0
9 Inverter~
13 662 1610 0 2 22
0 27 66
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3440 0 0
2
5.89816e-315 5.4889e-315
0
9 Inverter~
13 662 1509 0 2 22
0 47 55
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
6263 0 0
2
5.89816e-315 5.4902e-315
0
9 Inverter~
13 662 1535 0 2 22
0 46 56
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4900 0 0
2
5.89816e-315 5.49149e-315
0
9 Inverter~
13 662 1586 0 2 22
0 44 63
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
8783 0 0
2
5.89816e-315 5.49279e-315
0
9 Inverter~
13 662 1560 0 2 22
0 45 61
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3221 0 0
2
5.89816e-315 5.49408e-315
0
9 Inverter~
13 663 1458 0 2 22
0 49 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3215 0 0
2
5.89816e-315 5.49538e-315
0
9 Inverter~
13 663 1484 0 2 22
0 48 58
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
7903 0 0
2
5.89816e-315 5.49667e-315
0
9 Inverter~
13 663 1433 0 2 22
0 50 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
7121 0 0
2
5.89816e-315 5.49797e-315
0
9 Inverter~
13 663 1407 0 2 22
0 51 60
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4484 0 0
2
5.89816e-315 5.49926e-315
0
7 74LS154
95 551 1316 0 22 45
0 2 2 40 41 42 43 115 116 117
118 119 120 27 44 45 46 47 48 49
50 51 121
0
0 0 4848 270
6 74F154
-21 -87 21 -79
3 U17
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
5996 0 0
2
5.89816e-315 5.50056e-315
0
9 4-In NOR~
219 1422 275 0 5 22
0 70 69 68 67 29
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 1 0
1 U
7804 0 0
2
5.89816e-315 5.50185e-315
0
7 74LS126
116 1089 430 0 12 25
0 21 71 21 72 21 73 21 74 14
34 15 16
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
3 U15
-10 -52 11 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
5523 0 0
2
5.89816e-315 5.50315e-315
0
7 Ground~
168 1108 510 0 1 3
0 2
0
0 0 53360 270
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3330 0 0
2
5.89816e-315 0
0
7 74LS181
132 1190 471 0 22 45
0 75 22 76 75 67 68 69 70 80
79 78 77 23 2 122 123 124 125 71
72 73 74
0
0 0 4848 180
7 74LS181
-24 -69 25 -61
3 U14
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
3465 0 0
2
5.89816e-315 5.26354e-315
0
6 PROM32
80 777 600 0 14 29
0 6 2 33 32 31 30 38 37 36
35 14 34 15 16
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8396 0 0
2
5.89816e-315 5.30499e-315
0
AABKCADAEAFAGAHIICJAAFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 Ground~
168 389 599 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3685 0 0
2
5.89816e-315 5.32571e-315
0
7 74LS173
129 771 440 0 14 29
0 2 25 25 13 16 15 34 14 2
2 81 82 83 84
0
0 0 4848 270
6 74F173
-21 -51 21 -43
3 U12
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7849 0 0
2
5.89816e-315 5.34643e-315
0
7 Ground~
168 869 405 0 1 3
0 2
0
0 0 53360 90
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6343 0 0
2
5.89816e-315 5.3568e-315
0
7 Ground~
168 546 479 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7376 0 0
2
5.89816e-315 5.36716e-315
0
7 74LS257
147 614 517 0 14 29
0 85 81 86 82 87 83 88 84 89
2 30 31 32 33
0
0 0 4848 270
6 74F257
-21 -60 21 -52
3 U11
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9156 0 0
2
5.89816e-315 5.37752e-315
0
7 Ground~
168 475 168 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5776 0 0
2
5.89816e-315 5.38788e-315
0
2 +V
167 598 114 0 1 3
0 90
0
0 0 54256 0
2 5V
-8 -22 6 -14
3 V17
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7207 0 0
2
5.89816e-315 5.39306e-315
0
7 74LS193
137 663 168 0 14 29
0 17 90 7 2 14 34 15 16 126
127 94 93 92 91
0
0 0 4848 0
6 74F193
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4459 0 0
2
5.89816e-315 5.39824e-315
0
7 74LS126
116 833 168 0 12 25
0 9 94 9 93 9 92 9 91 14
34 15 16
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3760 0 0
2
5.89816e-315 5.40342e-315
0
7 74LS126
116 845 1176 0 12 25
0 24 99 24 100 24 101 24 102 16
15 34 14
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U8
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
754 0 0
2
5.89816e-315 5.4086e-315
0
7 Ground~
168 743 1174 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9767 0 0
2
5.89816e-315 5.41378e-315
0
7 74LS173
129 671 1128 0 14 29
0 2 5 5 13 16 15 34 14 2
2 99 100 101 102
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U7
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7978 0 0
2
5.89816e-315 5.41896e-315
0
7 74LS173
129 542 1127 0 14 29
0 28 5 5 13 35 36 37 38 2
2 43 42 41 40
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U6
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3142 0 0
2
5.89816e-315 5.42414e-315
0
14 Logic Display~
6 1390 1160 0 1 2
10 106
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
5.89816e-315 5.42933e-315
0
14 Logic Display~
6 1370 1160 0 1 2
10 105
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
659 0 0
2
5.89816e-315 5.43192e-315
0
14 Logic Display~
6 1350 1160 0 1 2
10 104
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
5.89816e-315 5.43451e-315
0
14 Logic Display~
6 1331 1160 0 1 2
10 103
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6792 0 0
2
5.89816e-315 5.4371e-315
0
7 Ground~
168 1253 1131 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3701 0 0
2
5.89816e-315 5.43969e-315
0
7 74LS173
129 1158 1090 0 14 29
0 2 4 4 13 14 34 15 16 2
2 103 104 105 106
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U5
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6316 0 0
2
5.89816e-315 5.44228e-315
0
7 Ground~
168 1400 746 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8734 0 0
2
5.89816e-315 5.44487e-315
0
7 74LS126
116 1090 852 0 12 25
0 20 95 20 96 20 97 20 98 14
34 15 16
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
7988 0 0
2
5.89816e-315 5.44746e-315
0
7 74LS257
147 1323 708 0 14 29
0 3 95 110 96 109 97 108 98 107
2 80 79 78 77
0
0 0 4848 90
6 74F257
-21 -60 21 -52
2 U3
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3217 0 0
2
5.89816e-315 5.45005e-315
0
7 74LS126
116 1091 294 0 12 25
0 18 67 18 68 18 69 18 70 14
34 15 16
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3965 0 0
2
5.89816e-315 5.45264e-315
0
7 Ground~
168 1254 242 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8239 0 0
2
5.89816e-315 5.45523e-315
0
7 74LS173
129 1159 200 0 14 29
0 2 19 19 13 14 34 15 16 2
2 67 68 69 70
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U1
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
828 0 0
2
5.89816e-315 5.45782e-315
0
14 Logic Display~
6 916 1239 0 1 2
10 38
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L16
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
42999.8 26
0
14 Logic Display~
6 935 1239 0 1 2
10 37
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L15
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7107 0 0
2
42999.8 27
0
14 Logic Display~
6 955 1239 0 1 2
10 36
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L14
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6433 0 0
2
42999.8 28
0
14 Logic Display~
6 975 1239 0 1 2
10 35
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L13
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8559 0 0
2
42999.8 29
0
14 Logic Display~
6 1053 1239 0 1 2
10 16
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L12
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3674 0 0
2
42999.8 30
0
14 Logic Display~
6 1033 1239 0 1 2
10 15
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L11
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5697 0 0
2
42999.8 31
0
14 Logic Display~
6 1013 1239 0 1 2
10 34
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L10
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
42999.8 32
0
14 Logic Display~
6 994 1239 0 1 2
10 14
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5219 0 0
2
42999.8 33
0
14 Logic Display~
6 994 94 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3795 0 0
2
42999.8 34
0
14 Logic Display~
6 1013 94 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3637 0 0
2
42999.8 35
0
14 Logic Display~
6 1033 94 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
42999.8 36
0
14 Logic Display~
6 1053 94 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6966 0 0
2
42999.8 37
0
14 Logic Display~
6 975 94 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9796 0 0
2
42999.8 38
0
14 Logic Display~
6 955 94 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
42999.8 39
0
14 Logic Display~
6 935 94 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
42999.8 40
0
14 Logic Display~
6 916 94 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
42999.8 41
0
289
1 0 3 0 0 0 0 15 0 0 62 2
1621 762
1621 762
1 0 4 0 0 4096 0 16 0 0 79 2
1577 1032
1577 1031
1 0 5 0 0 0 0 17 0 0 221 2
416 1075
416 1075
0 1 6 0 0 8320 0 0 91 24 0 4
920 1841
529 1841
529 564
739 564
0 2 7 0 0 8192 0 0 18 191 0 5
691 1752
691 1829
896 1829
896 1748
928 1748
0 2 8 0 0 8320 0 0 19 12 0 6
598 1694
598 1769
834 1769
834 1677
857 1677
857 1700
5 0 9 0 0 4096 0 100 0 0 10 4
801 177
790 177
790 178
787 178
3 0 9 0 0 0 0 100 0 0 10 4
801 159
790 159
790 160
787 160
1 0 9 0 0 0 0 100 0 0 10 4
801 141
790 141
790 142
787 142
0 7 9 0 0 8320 0 0 100 23 0 6
490 1632
17 1632
17 78
787 78
787 195
801 195
0 1 10 0 0 4096 0 0 20 104 0 3
848 1684
593 1684
593 1712
2 3 8 0 0 0 0 20 21 0 0 2
593 1694
603 1694
0 1 11 0 0 12288 0 0 21 102 0 6
946 1632
908 1632
908 1813
654 1813
654 1703
648 1703
0 2 12 0 0 4224 0 0 21 83 0 4
773 1738
665 1738
665 1685
648 1685
0 1 13 0 0 4096 0 0 22 234 0 4
1078 1020
1078 968
1088 968
1088 963
0 1 14 0 0 4096 0 0 23 242 0 4
1089 1036
1089 981
1114 981
1114 966
0 1 15 0 0 4096 0 0 24 244 0 4
1101 1050
1101 990
1139 990
1139 965
0 1 16 0 0 4096 0 0 25 245 0 4
1113 1060
1113 1008
1163 1008
1163 965
1 0 17 0 0 0 0 26 0 0 20 2
382 1857
382 1857
0 0 17 0 0 4096 0 0 0 222 0 2
382 1625
382 1862
0 1 17 0 0 0 0 0 27 107 0 2
462 1637
462 1865
1 0 9 0 0 0 0 28 0 0 23 2
488 1864
488 1864
3 0 9 0 0 0 0 20 0 0 0 5
547 1703
541 1703
541 1632
488 1632
488 1870
3 1 6 0 0 0 0 18 35 0 0 4
937 1793
937 1799
920 1799
920 1891
0 1 18 0 0 4096 0 0 34 263 0 2
1259 1712
1259 1913
0 1 19 0 0 4096 0 0 33 273 0 3
1301 1840
1301 1906
1300 1906
0 1 20 0 0 4096 0 0 32 204 0 2
1341 1835
1341 1904
0 1 21 0 0 4096 0 0 31 144 0 2
1367 1829
1367 1901
0 1 22 0 0 4096 0 0 30 259 0 2
1399 1824
1399 1894
0 1 23 0 0 4096 0 0 29 154 0 3
1430 1817
1430 1897
1431 1897
0 1 24 0 0 4096 0 0 36 212 0 3
632 1794
632 1872
633 1872
0 1 25 0 0 4096 0 0 37 82 0 2
822 1781
822 1858
1 0 7 0 0 0 0 38 0 0 34 2
667 1830
667 1830
0 0 7 0 0 0 0 0 0 191 0 2
667 1752
667 1834
3 3 26 0 0 12416 0 39 67 0 0 6
358 1200
380 1200
380 1224
659 1224
659 1324
684 1324
1 0 27 0 0 4096 0 39 0 0 37 2
313 1191
267 1191
0 0 27 0 0 8320 0 0 0 67 0 3
562 1599
267 1599
267 1176
0 2 13 0 0 4096 0 0 39 39 0 2
169 1209
313 1209
0 0 13 0 0 8192 0 0 0 234 84 3
167 1020
169 1020
169 1230
2 0 10 0 0 4096 0 40 0 0 121 3
398 1388
776 1388
776 1355
3 1 28 0 0 8320 0 40 104 0 0 5
389 1339
389 1201
610 1201
610 1097
571 1097
1 1 2 0 0 4096 0 40 41 0 0 2
380 1388
380 1386
9 0 2 0 0 4096 0 104 0 0 229 2
571 1167
571 1175
0 0 5 0 0 4096 0 0 0 61 221 3
554 1065
469 1065
469 1075
1 0 2 0 0 0 0 42 0 0 132 2
571 1271
571 1272
1 5 29 0 0 12416 0 60 87 0 0 5
791 1639
791 1260
1486 1260
1486 275
1461 275
6 11 30 0 0 4224 0 91 96 0 0 3
745 636
631 636
631 554
5 12 31 0 0 4224 0 91 96 0 0 3
745 627
613 627
613 554
13 4 32 0 0 8320 0 96 91 0 0 3
595 554
595 618
745 618
14 3 33 0 0 8320 0 96 91 0 0 3
577 554
577 609
745 609
0 14 16 0 0 4096 0 0 91 282 0 2
1053 636
809 636
0 13 15 0 0 4096 0 0 91 283 0 2
1033 627
809 627
0 12 34 0 0 4096 0 0 91 284 0 2
1013 618
809 618
0 11 14 0 0 4096 0 0 91 285 0 2
994 609
809 609
0 10 35 0 0 4096 0 0 91 286 0 2
975 600
809 600
0 9 36 0 0 4096 0 0 91 287 0 2
955 591
809 591
0 8 37 0 0 4096 0 0 91 288 0 2
935 582
809 582
0 7 38 0 0 4096 0 0 91 289 0 2
916 573
809 573
1 2 2 0 0 4224 0 92 91 0 0 2
396 600
745 600
1 3 39 0 0 4224 0 18 44 0 0 3
946 1748
946 1747
945 1747
3 2 5 0 0 0 0 104 104 0 0 5
553 1091
554 1091
554 1065
562 1065
562 1091
2 1 3 0 0 4224 0 43 113 0 0 3
1761 762
1282 762
1282 739
14 3 40 0 0 4224 0 104 86 0 0 4
508 1161
508 1257
535 1257
535 1286
13 4 41 0 0 4224 0 104 86 0 0 4
517 1161
517 1262
526 1262
526 1286
12 5 42 0 0 4224 0 104 86 0 0 4
526 1161
526 1267
517 1267
517 1286
11 6 43 0 0 4224 0 104 86 0 0 4
535 1161
535 1272
508 1272
508 1286
13 1 27 0 0 0 0 86 77 0 0 3
562 1356
562 1610
647 1610
14 1 44 0 0 4224 0 86 80 0 0 3
553 1356
553 1586
647 1586
15 1 45 0 0 4224 0 86 81 0 0 3
544 1356
544 1560
647 1560
16 1 46 0 0 4224 0 86 79 0 0 3
535 1356
535 1535
647 1535
17 1 47 0 0 4224 0 86 78 0 0 3
526 1356
526 1509
647 1509
18 1 48 0 0 8320 0 86 83 0 0 3
517 1356
517 1484
648 1484
19 1 49 0 0 8320 0 86 82 0 0 3
508 1356
508 1458
648 1458
20 1 50 0 0 8320 0 86 84 0 0 3
499 1356
499 1433
648 1433
21 1 51 0 0 8320 0 86 85 0 0 3
490 1356
490 1407
648 1407
2 3 52 0 0 4224 0 46 57 0 0 3
987 1799
987 1689
955 1689
3 1 52 0 0 0 0 57 44 0 0 4
955 1689
955 1694
954 1694
954 1695
1 0 2 0 0 0 0 110 0 0 240 3
1187 1060
1225 1060
1225 1132
2 3 4 0 0 4224 0 45 110 0 0 3
1684 1031
1169 1031
1169 1054
0 1 18 0 0 4096 0 0 45 263 0 3
1950 1033
1720 1033
1720 1031
1 0 24 0 0 0 0 19 0 0 212 4
866 1699
866 1698
875 1698
875 1685
4 2 25 0 0 12416 0 19 93 0 0 6
857 1751
857 1781
14 1781
14 295
791 295
791 404
3 2 12 0 0 0 0 59 48 0 0 3
773 1732
773 1743
764 1743
0 1 13 0 0 16384 0 0 2 0 0 5
167 1225
169 1225
169 1230
322 1230
322 1449
1 0 23 0 0 0 0 49 0 0 154 2
1875 587
1875 634
0 1 22 0 0 4096 0 0 50 259 0 3
1934 764
1934 545
1873 545
4 2 53 0 0 8320 0 55 51 0 0 3
1032 1670
1084 1670
1084 1765
1 0 54 0 0 4096 0 51 0 0 119 2
1102 1765
1102 1304
1 0 55 0 0 4096 0 52 0 0 126 2
1192 1722
1192 1511
2 0 54 0 0 0 0 52 0 0 119 2
1174 1722
1174 1304
1 0 54 0 0 0 0 53 0 0 119 2
1134 1667
1134 1304
2 0 56 0 0 4096 0 53 0 0 125 2
1116 1667
1116 1537
1 0 55 0 0 0 0 54 0 0 126 2
1051 1680
1051 1511
3 1 57 0 0 4224 0 54 56 0 0 4
1042 1726
1042 1742
1033 1742
1033 1743
2 4 53 0 0 0 0 54 55 0 0 3
1033 1680
1033 1670
1032 1670
1 0 58 0 0 4096 0 55 0 0 127 2
1041 1624
1041 1486
2 0 22 0 0 0 0 55 0 0 128 2
1032 1625
1032 1460
3 0 23 0 0 4096 0 55 0 0 129 2
1023 1624
1023 1435
2 0 54 0 0 0 0 56 0 0 119 2
1015 1743
1015 1304
3 1 59 0 0 8320 0 56 46 0 0 4
1024 1788
1024 1796
1005 1796
1005 1799
2 0 17 0 0 4096 0 44 0 0 120 4
936 1695
936 1344
937 1344
937 1329
2 0 11 0 0 4096 0 57 0 0 118 2
946 1644
946 1278
1 0 60 0 0 4096 0 57 0 0 130 2
964 1644
964 1409
3 0 10 0 0 0 0 19 0 0 121 4
848 1699
848 1370
857 1370
857 1355
1 0 54 0 0 0 0 58 0 0 119 2
884 1640
884 1304
2 0 60 0 0 0 0 58 0 0 130 2
866 1640
866 1409
0 1 17 0 0 12416 0 0 99 120 0 7
825 1329
825 1637
6 1637
6 110
385 110
385 141
631 141
1 0 54 0 0 0 0 48 0 0 119 5
764 1761
791 1761
791 1730
820 1730
820 1304
2 0 61 0 0 4096 0 59 0 0 124 2
764 1686
764 1562
1 3 62 0 0 4224 0 59 60 0 0 2
782 1686
782 1684
2 0 63 0 0 4096 0 60 0 0 123 2
773 1639
773 1588
1 4 64 0 0 8320 0 61 67 0 0 3
675 1357
678 1357
678 1342
3 0 54 0 0 0 0 62 0 0 119 3
736 1252
779 1252
779 1304
2 0 17 0 0 0 0 62 0 0 120 3
735 1261
774 1261
774 1329
1 0 10 0 0 0 0 62 0 0 121 3
736 1270
770 1270
770 1355
2 0 65 0 0 4096 0 67 0 0 117 3
684 1306
669 1306
669 1297
1 4 65 0 0 8320 0 67 62 0 0 4
684 1297
669 1297
669 1261
684 1261
9 1 11 0 0 12416 0 67 66 0 0 4
748 1333
766 1333
766 1278
1536 1278
10 1 54 0 0 12416 0 67 63 0 0 4
748 1342
759 1342
759 1304
1536 1304
1 11 17 0 0 0 0 64 67 0 0 4
1536 1329
754 1329
754 1351
748 1351
1 12 10 0 0 4224 0 65 67 0 0 4
1536 1355
754 1355
754 1360
748 1360
2 1 66 0 0 8320 0 77 75 0 0 3
683 1610
683 1612
1534 1612
2 1 63 0 0 8320 0 80 72 0 0 3
683 1586
683 1588
1534 1588
2 1 61 0 0 8320 0 81 71 0 0 3
683 1560
683 1562
1533 1562
2 1 56 0 0 8320 0 79 73 0 0 3
683 1535
683 1537
1533 1537
2 1 55 0 0 8320 0 78 74 0 0 3
683 1509
683 1511
1533 1511
2 1 58 0 0 8320 0 83 69 0 0 3
684 1484
684 1486
1534 1486
2 1 22 0 0 8192 0 82 70 0 0 3
684 1458
684 1460
1534 1460
2 1 23 0 0 8192 0 84 76 0 0 3
684 1433
684 1435
1534 1435
2 1 60 0 0 8320 0 85 68 0 0 3
684 1407
684 1409
1534 1409
0 2 66 0 0 0 0 0 77 0 0 4
684 1610
682 1610
682 1610
683 1610
1 2 2 0 0 0 0 86 86 0 0 4
571 1280
571 1272
562 1272
562 1280
0 4 67 0 0 4096 0 0 87 140 0 4
1233 316
1356 316
1356 289
1405 289
0 3 68 0 0 4096 0 0 87 139 0 4
1245 299
1343 299
1343 280
1405 280
0 2 69 0 0 4096 0 0 87 138 0 4
1255 282
1334 282
1334 271
1405 271
0 1 70 0 0 4096 0 0 87 137 0 2
1265 262
1405 262
8 8 70 0 0 8320 0 90 114 0 0 4
1228 457
1265 457
1265 262
1123 262
7 0 69 0 0 8320 0 90 0 0 270 4
1228 466
1255 466
1255 280
1134 280
6 0 68 0 0 8320 0 90 0 0 269 4
1228 475
1245 475
1245 298
1143 298
0 5 67 0 0 8320 0 0 90 268 0 4
1152 316
1236 316
1236 484
1228 484
7 0 21 0 0 0 0 88 0 0 144 2
1121 407
1128 407
5 0 21 0 0 0 0 88 0 0 144 2
1121 425
1128 425
3 0 21 0 0 0 0 88 0 0 144 2
1121 443
1128 443
3 1 21 0 0 12416 0 51 88 0 0 7
1093 1810
1093 1829
1939 1829
1939 375
1128 375
1128 461
1121 461
2 19 71 0 0 4224 0 88 90 0 0 3
1121 452
1152 452
1152 448
4 20 72 0 0 4224 0 88 90 0 0 4
1121 434
1147 434
1147 439
1152 439
6 21 73 0 0 4224 0 88 90 0 0 4
1121 416
1142 416
1142 430
1152 430
22 8 74 0 0 12416 0 90 88 0 0 4
1152 421
1146 421
1146 398
1121 398
9 0 14 0 0 0 0 88 0 0 285 2
1057 452
994 452
10 0 34 0 0 0 0 88 0 0 284 2
1057 434
1013 434
11 0 15 0 0 0 0 88 0 0 283 2
1057 416
1033 416
12 0 16 0 0 0 0 88 0 0 282 2
1057 398
1053 398
14 1 2 0 0 0 0 90 89 0 0 2
1158 511
1115 511
13 0 23 0 0 16512 0 90 0 0 129 7
1158 520
1146 520
1146 634
1929 634
1929 1817
1231 1817
1231 1435
4 2 75 0 0 4224 0 90 50 0 0 4
1222 493
1839 493
1839 545
1837 545
3 2 76 0 0 4224 0 90 49 0 0 4
1222 502
1807 502
1807 587
1839 587
2 0 22 0 0 0 0 90 0 0 86 4
1222 511
1776 511
1776 561
1934 561
1 2 75 0 0 0 0 90 50 0 0 4
1222 520
1743 520
1743 545
1837 545
12 14 77 0 0 8320 0 90 113 0 0 3
1228 421
1354 421
1354 675
11 13 78 0 0 8320 0 90 113 0 0 3
1228 430
1336 430
1336 675
10 12 79 0 0 8320 0 90 113 0 0 3
1228 439
1318 439
1318 675
9 11 80 0 0 8320 0 90 113 0 0 3
1228 448
1300 448
1300 675
8 0 38 0 0 8192 0 104 0 0 289 3
508 1097
508 935
916 935
0 7 37 0 0 4096 0 0 104 288 0 3
935 946
517 946
517 1097
6 0 36 0 0 8192 0 104 0 0 287 3
526 1097
526 961
955 961
5 0 35 0 0 8192 0 104 0 0 286 3
535 1097
535 975
975 975
2 11 81 0 0 8320 0 96 93 0 0 4
640 490
640 483
764 483
764 474
12 4 82 0 0 8320 0 93 96 0 0 4
755 474
755 480
622 480
622 490
6 13 83 0 0 8320 0 96 93 0 0 4
604 490
604 477
746 477
746 474
14 8 84 0 0 4224 0 93 96 0 0 3
737 474
586 474
586 490
4 0 13 0 0 8192 0 93 0 0 234 3
773 410
773 275
167 275
5 0 16 0 0 8192 0 93 0 0 282 3
764 410
764 363
1053 363
6 0 15 0 0 8192 0 93 0 0 283 3
755 410
755 353
1033 353
7 0 34 0 0 8192 0 93 0 0 284 3
746 410
746 342
1013 342
8 0 14 0 0 8192 0 93 0 0 285 3
737 410
737 330
994 330
3 0 25 0 0 0 0 93 0 0 82 3
782 404
782 395
791 395
9 0 2 0 0 0 0 93 0 0 178 2
800 480
800 490
10 0 2 0 0 0 0 93 0 0 179 4
791 480
791 490
851 490
851 406
1 1 2 0 0 0 0 93 94 0 0 3
800 410
800 406
862 406
1 10 2 0 0 0 0 95 96 0 0 3
553 480
568 480
568 484
1 1 85 0 0 8320 0 96 1 0 0 5
649 490
649 359
263 359
263 441
218 441
1 3 86 0 0 8320 0 3 96 0 0 4
381 488
381 412
631 412
631 490
1 5 87 0 0 8320 0 4 96 0 0 4
349 487
349 397
613 397
613 490
1 7 88 0 0 8320 0 5 96 0 0 4
318 487
318 383
595 383
595 490
1 9 89 0 0 8320 0 6 96 0 0 4
285 485
285 370
577 370
577 490
9 0 14 0 0 0 0 100 0 0 285 4
865 150
979 150
979 151
994 151
10 0 34 0 0 0 0 100 0 0 284 4
865 168
998 168
998 169
1013 169
11 0 15 0 0 0 0 100 0 0 283 4
865 186
1018 186
1018 187
1033 187
12 0 16 0 0 0 0 100 0 0 282 4
865 204
1038 204
1038 205
1053 205
1 4 2 0 0 0 0 97 99 0 0 3
482 169
482 168
631 168
3 3 7 0 0 12416 0 99 48 0 0 7
625 159
625 158
2 158
2 1775
616 1775
616 1752
713 1752
2 1 90 0 0 4224 0 99 98 0 0 3
631 150
598 150
598 123
0 5 14 0 0 4096 0 0 99 285 0 4
994 248
593 248
593 177
631 177
0 6 34 0 0 4096 0 0 99 284 0 4
1013 240
602 240
602 186
631 186
0 7 15 0 0 4096 0 0 99 283 0 4
1033 231
611 231
611 195
631 195
0 8 16 0 0 4096 0 0 99 282 0 4
1053 222
620 222
620 204
631 204
8 14 91 0 0 4224 0 100 99 0 0 2
801 204
695 204
6 13 92 0 0 4224 0 100 99 0 0 4
801 186
748 186
748 195
695 195
4 12 93 0 0 4224 0 100 99 0 0 4
801 168
740 168
740 186
695 186
11 2 94 0 0 12416 0 99 100 0 0 4
695 177
731 177
731 150
801 150
7 0 20 0 0 0 0 112 0 0 204 2
1122 829
1148 829
5 0 20 0 0 0 0 112 0 0 204 2
1122 847
1148 847
3 0 20 0 0 0 0 112 0 0 204 2
1122 865
1148 865
3 1 20 0 0 12416 0 52 112 0 0 7
1183 1767
1183 1835
1945 1835
1945 802
1148 802
1148 883
1122 883
2 0 95 0 0 4096 0 112 0 0 258 2
1122 874
1290 874
4 0 96 0 0 4096 0 112 0 0 257 2
1122 856
1309 856
6 0 97 0 0 4224 0 112 0 0 256 2
1122 838
1327 838
8 0 98 0 0 4224 0 112 0 0 255 2
1122 820
1345 820
7 0 24 0 0 0 0 101 0 0 212 2
813 1203
758 1203
5 0 24 0 0 0 0 101 0 0 212 3
813 1185
813 1171
758 1171
3 0 24 0 0 0 0 101 0 0 212 2
813 1167
758 1167
3 1 24 0 0 12416 0 58 101 0 0 8
875 1685
886 1685
886 1794
26 1794
26 1238
758 1238
758 1149
813 1149
11 2 99 0 0 8320 0 103 101 0 0 5
664 1162
664 1186
793 1186
793 1158
813 1158
12 0 14 0 0 0 0 101 0 0 285 2
877 1212
994 1212
11 0 34 0 0 0 0 101 0 0 284 2
877 1194
1013 1194
10 0 15 0 0 0 0 101 0 0 283 2
877 1176
1033 1176
9 0 16 0 0 0 0 101 0 0 282 2
877 1158
1053 1158
12 4 100 0 0 8320 0 103 101 0 0 5
655 1162
655 1190
807 1190
807 1176
813 1176
13 6 101 0 0 8320 0 103 101 0 0 3
646 1162
646 1194
813 1194
14 8 102 0 0 8320 0 103 101 0 0 3
637 1162
637 1212
813 1212
3 2 5 0 0 8320 0 103 47 0 0 5
682 1092
682 1075
346 1075
346 1059
341 1059
0 1 17 0 0 0 0 0 47 120 0 5
837 1329
837 1625
22 1625
22 1059
305 1059
3 2 5 0 0 0 0 103 103 0 0 2
682 1092
691 1092
0 0 13 0 0 0 0 0 0 225 234 2
673 1087
673 1020
4 4 13 0 0 0 0 103 104 0 0 4
673 1098
673 1085
544 1085
544 1097
1 0 2 0 0 0 0 102 0 0 227 4
736 1175
737 1175
737 1175
736 1175
1 0 2 0 0 0 0 103 0 0 228 4
700 1098
736 1098
736 1175
699 1175
0 9 2 0 0 0 0 0 103 229 0 3
690 1175
700 1175
700 1168
10 10 2 0 0 0 0 104 103 0 0 4
562 1167
562 1175
691 1175
691 1168
5 0 16 0 0 0 0 103 0 0 282 3
664 1098
664 1068
1053 1068
6 0 15 0 0 0 0 103 0 0 283 3
655 1098
655 1063
1033 1063
7 0 34 0 0 0 0 103 0 0 284 3
646 1098
646 1057
1013 1057
8 0 14 0 0 0 0 103 0 0 285 3
637 1098
637 1051
994 1051
4 0 13 0 0 8192 0 110 0 0 277 4
1160 1060
1160 1020
167 1020
167 31
11 1 103 0 0 8320 0 110 108 0 0 4
1151 1124
1151 1217
1331 1217
1331 1178
12 1 104 0 0 8320 0 110 107 0 0 4
1142 1124
1142 1210
1350 1210
1350 1178
13 1 105 0 0 8320 0 110 106 0 0 4
1133 1124
1133 1199
1370 1199
1370 1178
14 1 106 0 0 8320 0 110 105 0 0 4
1124 1124
1124 1189
1390 1189
1390 1178
9 0 2 0 0 0 0 110 0 0 240 2
1187 1130
1187 1132
10 1 2 0 0 0 0 110 109 0 0 3
1178 1130
1178 1132
1246 1132
2 0 4 0 0 0 0 110 0 0 79 2
1178 1054
1178 1031
5 0 14 0 0 0 0 110 0 0 285 3
1151 1060
1151 1036
994 1036
6 0 34 0 0 0 0 110 0 0 284 3
1142 1060
1142 1042
1013 1042
7 0 15 0 0 0 0 110 0 0 283 3
1133 1060
1133 1050
1033 1050
8 0 16 0 0 0 0 110 0 0 282 2
1124 1060
1053 1060
1 10 2 0 0 0 0 111 113 0 0 3
1393 747
1393 745
1363 745
9 0 14 0 0 0 0 112 0 0 285 2
1058 874
994 874
10 0 34 0 0 0 0 112 0 0 284 2
1058 856
1013 856
11 0 15 0 0 0 0 112 0 0 283 2
1058 838
1033 838
12 0 16 0 0 0 0 112 0 0 282 2
1058 820
1053 820
9 1 107 0 0 8320 0 113 10 0 0 4
1354 739
1354 835
1633 835
1633 955
7 1 108 0 0 8320 0 113 9 0 0 4
1336 739
1336 849
1601 849
1601 954
5 1 109 0 0 8320 0 113 8 0 0 4
1318 739
1318 864
1570 864
1570 954
3 1 110 0 0 8320 0 113 7 0 0 4
1300 739
1300 878
1537 878
1537 952
8 1 98 0 0 0 0 113 11 0 0 4
1345 739
1345 918
1386 918
1386 953
6 1 97 0 0 0 0 113 12 0 0 4
1327 739
1327 928
1354 928
1354 952
4 1 96 0 0 4224 0 113 13 0 0 4
1309 739
1309 938
1323 938
1323 952
2 1 95 0 0 8320 0 113 14 0 0 3
1291 739
1290 739
1290 950
0 1 22 0 0 12416 0 0 43 128 0 5
1222 1460
1222 1824
1934 1824
1934 762
1797 762
0 7 18 0 0 0 0 0 114 261 0 3
1129 290
1129 271
1123 271
0 5 18 0 0 0 0 0 114 262 0 3
1129 307
1129 289
1123 289
3 0 18 0 0 0 0 114 0 0 263 3
1123 307
1129 307
1129 325
1 3 18 0 0 8320 0 114 53 0 0 4
1123 325
1950 325
1950 1712
1125 1712
9 0 14 0 0 0 0 114 0 0 285 2
1059 316
994 316
10 0 34 0 0 0 0 114 0 0 284 2
1059 298
1013 298
11 0 15 0 0 0 0 114 0 0 283 2
1059 280
1033 280
12 0 16 0 0 0 0 114 0 0 282 2
1059 262
1053 262
11 2 67 0 0 0 0 116 114 0 0 3
1152 234
1152 316
1123 316
12 4 68 0 0 0 0 116 114 0 0 3
1143 234
1143 298
1123 298
13 6 69 0 0 0 0 116 114 0 0 3
1134 234
1134 280
1123 280
14 8 70 0 0 0 0 116 114 0 0 3
1125 234
1123 234
1123 262
2 0 19 0 0 0 0 116 0 0 273 2
1179 164
1179 141
3 3 19 0 0 16512 0 46 116 0 0 7
996 1851
1016 1851
1016 1840
1955 1840
1955 141
1170 141
1170 164
1 0 2 0 0 0 0 116 0 0 276 3
1188 170
1220 170
1220 243
9 0 2 0 0 0 0 116 0 0 276 2
1188 240
1188 243
10 1 2 0 0 0 0 116 115 0 0 3
1179 240
1179 243
1247 243
0 4 13 0 0 4224 0 0 116 0 0 3
112 31
1161 31
1161 170
5 0 14 0 0 0 0 116 0 0 285 3
1152 170
1152 146
994 146
6 0 34 0 0 0 0 116 0 0 284 3
1143 170
1143 152
1013 152
7 0 15 0 0 0 0 116 0 0 283 3
1134 170
1134 160
1033 160
8 0 16 0 0 0 0 116 0 0 282 2
1125 170
1053 170
1 1 16 0 0 4224 0 128 121 0 0 2
1053 112
1053 1225
1 1 15 0 0 4224 0 127 122 0 0 2
1033 112
1033 1225
1 1 34 0 0 4224 0 126 123 0 0 2
1013 112
1013 1225
1 1 14 0 0 4224 0 125 124 0 0 2
994 112
994 1225
1 1 35 0 0 4224 0 129 120 0 0 2
975 112
975 1225
1 1 36 0 0 4224 0 130 119 0 0 2
955 112
955 1225
1 1 37 0 0 4224 0 131 118 0 0 2
935 112
935 1225
1 1 38 0 0 4224 0 132 117 0 0 2
916 112
916 1225
60
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 9
158 445 294 476
170 455 281 476
9 SM(MAR=1)
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
707 1583 775 1614
720 1593 761 1614
3 HLT
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
712 1559 763 1590
725 1569 749 1590
2 JZ
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
707 1530 772 1561
719 1540 759 1561
3 JMP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
706 1504 772 1535
718 1514 759 1535
3 OUT
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
707 1428 773 1459
720 1438 759 1459
3 SUB
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
706 1402 774 1433
718 1412 761 1433
3 ADD
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
709 1379 774 1410
721 1389 761 1410
3 LDA
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
781 1323 829 1351
794 1333 815 1353
2 T1
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
782 1297 831 1325
794 1307 818 1327
2 T2
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
783 1272 834 1300
796 1282 820 1302
2 T3
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
786 1248 837 1276
799 1258 823 1278
2 T4
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1628 105 1676 136
1639 114 1664 135
2 LA
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1648 293 1685 324
1653 297 1679 318
2 EA
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1747 771 1792 802
1755 778 1783 799
2 EB
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1749 1032 1798 1063
1759 1040 1787 1061
2 LO
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
123 41 170 72
133 49 159 70
2 EP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
121 125 167 156
131 133 156 154
2 LP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
784 665 829 696
793 672 819 693
2 CE
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
706 78 766 123
715 85 756 116
2 PC
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
798 285 887 330
807 292 877 323
3 MAR
-24 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 11
354 315 567 360
363 322 557 353
11 INPUT & MUX
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
641 977 698 1022
650 985 688 1016
2 IR
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
117 262 168 293
127 269 157 290
2 LM
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
102 1054 142 1085
111 1061 132 1082
2 LI
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
115 1237 157 1268
124 1245 147 1266
2 EI
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 5
112 -2 199 29
121 6 189 27
5 CLOCK
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
122 86 166 117
131 93 156 114
2 CP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
1704 635 1751 666
1713 642 1741 663
3 Cin
-19 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1736 510 1783 547
1745 517 1773 542
2 S2
-19 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1770 503 1813 540
1779 511 1803 536
2 S1
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1802 501 1845 532
1811 508 1835 529
2 S0
-19 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1692 525 1739 562
1701 533 1729 558
2 S3
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1642 338 1687 369
1652 345 1676 366
2 Eu
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1272 190 1312 235
1282 197 1301 228
1 A
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1248 901 1290 946
1257 908 1280 939
1 B
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1646 894 1685 939
1655 901 1675 932
1 C
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 7
1191 982 1350 1027
1200 989 1340 1020
7 OUT REG
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 7
1300 1090 1455 1135
1309 1097 1445 1128
7 DISPLAY
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 5
164 1294 257 1325
176 1304 244 1325
5 CLOCK
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
1175 671 1265 716
1185 681 1254 712
3 MUX
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
1382 419 1474 464
1397 429 1458 460
3 ALU
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 14
283 1482 514 1527
298 1492 498 1523
14 Control Matrix
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
709 1455 773 1486
719 1464 762 1485
3 AND
-19 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
705 1474 771 1511
718 1484 757 1509
3 mov
-21 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1695 723 1726 765
1705 733 1715 761
1 s
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
471 1883 518 1914
481 1891 507 1912
2 EP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
424 1896 468 1927
433 1903 458 1924
2 CP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
661 1862 707 1893
671 1870 696 1891
2 LP
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
796 1890 847 1921
806 1897 836 1918
2 LM
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
371 1900 411 1931
380 1907 401 1928
2 LI
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
604 1904 646 1935
613 1912 636 1933
2 EI
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1239 1945 1276 1976
1244 1949 1270 1970
2 EA
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1349 1930 1394 1961
1359 1937 1383 1958
2 Eu
-21 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1386 1922 1417 1964
1396 1932 1406 1960
1 s
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1314 1936 1359 1967
1322 1943 1350 1964
2 EB
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
1419 1934 1466 1965
1428 1941 1456 1962
3 Cin
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1276 1944 1324 1975
1287 1953 1312 1974
2 LA
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
903 1925 948 1956
912 1932 938 1953
2 CE
-24 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 3
727 491 835 536
744 503 817 534
3 ROM
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
