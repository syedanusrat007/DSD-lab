CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1170 15 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
122
13 Logic Switch~
5 206 441 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3965 0 0
2
43001.6 0
0
13 Logic Switch~
5 168 1409 0 1 11
0 3
0
0 0 21360 90
2 0V
11 0 25 8
3 V31
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8239 0 0
2
5.89815e-315 5.26354e-315
0
13 Logic Switch~
5 380 501 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V20
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
828 0 0
2
5.89815e-315 5.30499e-315
0
13 Logic Switch~
5 348 500 0 1 11
0 85
0
0 0 21360 90
2 0V
11 0 25 8
3 V22
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6187 0 0
2
5.89815e-315 5.32571e-315
0
13 Logic Switch~
5 317 500 0 1 11
0 86
0
0 0 21360 90
2 0V
11 0 25 8
3 V23
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7107 0 0
2
5.89815e-315 5.34643e-315
0
13 Logic Switch~
5 284 498 0 1 11
0 87
0
0 0 21360 90
2 0V
11 0 25 8
3 V24
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6433 0 0
2
5.89815e-315 5.3568e-315
0
13 Logic Switch~
5 1536 965 0 1 11
0 108
0
0 0 21360 90
2 0V
11 0 25 8
3 V12
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8559 0 0
2
5.89815e-315 5.36716e-315
0
13 Logic Switch~
5 1569 967 0 1 11
0 107
0
0 0 21360 90
2 0V
11 0 25 8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3674 0 0
2
5.89815e-315 5.37752e-315
0
13 Logic Switch~
5 1600 967 0 1 11
0 106
0
0 0 21360 90
2 0V
11 0 25 8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5697 0 0
2
5.89815e-315 5.38788e-315
0
13 Logic Switch~
5 1632 968 0 10 11
0 105 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3805 0 0
2
5.89815e-315 5.39306e-315
0
13 Logic Switch~
5 1385 966 0 10 11
0 96 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5219 0 0
2
5.89815e-315 5.39824e-315
0
13 Logic Switch~
5 1353 965 0 1 11
0 95
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3795 0 0
2
5.89815e-315 5.40342e-315
0
13 Logic Switch~
5 1322 965 0 1 11
0 94
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3637 0 0
2
5.89815e-315 5.4086e-315
0
13 Logic Switch~
5 1289 963 0 1 11
0 93
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3226 0 0
2
5.89815e-315 5.41378e-315
0
14 Logic Display~
6 74 1983 0 1 2
10 15
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L46
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6966 0 0
2
43001.6 0
0
14 Logic Display~
6 174 1976 0 1 2
10 15
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L45
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9796 0 0
2
43001.6 0
0
14 Logic Display~
6 1281 1961 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L44
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5952 0 0
2
43001.6 0
0
14 Logic Display~
6 1156 1964 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L43
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3649 0 0
2
43001.6 0
0
14 Logic Display~
6 1024 1961 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L42
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3716 0 0
2
43001.6 0
0
14 Logic Display~
6 899 1959 0 1 2
10 8
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L41
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4797 0 0
2
43001.6 0
0
14 Logic Display~
6 776 1967 0 1 2
10 9
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4681 0 0
2
43001.6 0
0
14 Logic Display~
6 660 1974 0 1 2
10 10
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L39
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9730 0 0
2
43001.6 0
0
14 Logic Display~
6 560 1976 0 1 2
10 11
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L38
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9874 0 0
2
43001.6 0
0
14 Logic Display~
6 473 1974 0 1 2
10 12
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L37
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
364 0 0
2
43001.6 0
0
14 Logic Display~
6 384 1977 0 1 2
10 13
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L36
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3656 0 0
2
43001.6 0
0
14 Logic Display~
6 289 1977 0 1 2
10 14
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L35
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3131 0 0
2
43001.6 0
0
9 2-In AND~
219 337 1200 0 3 22
0 16 3 4
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U30B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
6772 0 0
2
43001.6 1
0
9 2-In XOR~
219 386 1369 0 3 22
0 2 14 17
0
0 0 624 90
6 74LS86
-21 -24 21 -16
4 U31A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
9557 0 0
2
5.89815e-315 5.41896e-315
0
7 Ground~
168 380 1392 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5789 0 0
2
5.89815e-315 5.42414e-315
0
7 Ground~
168 571 1263 0 1 3
0 2
0
0 0 53360 180
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7328 0 0
2
5.89815e-315 5.42933e-315
0
9 2-In AND~
219 939 1767 0 3 22
0 32 12 10
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U30A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
4799 0 0
2
43001.6 2
0
9 Inverter~
13 1776 762 0 2 22
0 49 33
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U29C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
9196 0 0
2
43001.6 3
0
9 2-In NOR~
219 939 1714 0 3 22
0 46 15 32
0
0 0 624 270
4 7428
-14 -24 14 -16
4 U28C
32 -10 60 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
3857 0 0
2
43001.6 4
0
9 Inverter~
13 1699 1031 0 2 22
0 9 5
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U29B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
7125 0 0
2
5.89815e-315 5.43192e-315
0
9 2-In NOR~
219 990 1818 0 3 22
0 56 46 8
0
0 0 624 270
4 7428
-14 -24 14 -16
4 U28B
32 -10 60 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3641 0 0
2
5.89815e-315 5.43451e-315
0
9 Inverter~
13 320 1059 0 2 22
0 15 18
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U29A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
9821 0 0
2
5.89815e-315 5.4371e-315
0
9 2-In NOR~
219 851 1719 0 3 22
0 13 14 11
0
0 0 624 270
4 7428
-14 -24 14 -16
4 U28A
32 -10 60 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3187 0 0
2
5.89815e-315 5.43969e-315
0
5 4011~
219 740 1752 0 3 22
0 51 47 12
0
0 0 624 180
4 4011
-7 -24 21 -16
4 U27A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 10 0
1 U
762 0 0
2
5.89815e-315 5.44228e-315
0
9 Inverter~
13 1854 587 0 2 22
0 48 74
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U19F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
39 0 0
2
43001.6 7
0
9 Inverter~
13 1852 545 0 2 22
0 49 73
0
0 0 624 180
5 74F04
-18 -19 17 -11
4 U19E
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
9450 0 0
2
43001.6 8
0
9 2-In AND~
219 1095 1787 0 3 22
0 51 50 6
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3236 0 0
2
43001.6 9
0
9 2-In AND~
219 1185 1744 0 3 22
0 52 51 7
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3321 0 0
2
43001.6 10
0
9 2-In AND~
219 1127 1689 0 3 22
0 51 53 9
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8879 0 0
2
43001.6 11
0
8 2-In OR~
219 1039 1696 0 3 22
0 52 50 54
0
0 0 624 270
5 74F32
-18 -24 17 -16
4 U26A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5433 0 0
2
43001.6 12
0
8 3-In OR~
219 1029 1640 0 4 22
0 55 49 48 50
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U25A
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
3679 0 0
2
43001.6 13
0
9 2-In AND~
219 1026 1765 0 3 22
0 54 51 56
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U24A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9342 0 0
2
43001.6 14
0
9 2-In AND~
219 957 1666 0 3 22
0 58 57 46
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3623 0 0
2
43001.6 15
0
9 2-In AND~
219 877 1662 0 3 22
0 51 58 13
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3722 0 0
2
43001.6 16
0
8 2-In OR~
219 770 1702 0 3 22
0 60 59 47
0
0 0 624 270
5 74F32
-18 -24 17 -16
4 U23A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8993 0 0
2
43001.6 17
0
9 2-In AND~
219 784 1661 0 3 22
0 19 61 60
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3723 0 0
2
43001.6 18
0
2 +V
167 675 1372 0 1 3
0 62
0
0 0 54256 180
3 10V
6 -2 27 6
3 V32
6 -12 27 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6244 0 0
2
43001.6 19
0
9 3-In NOR~
219 711 1261 0 4 22
0 14 15 51 63
0
0 0 624 180
5 74F27
-18 -24 17 -16
4 U21A
-11 -2 17 6
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
6421 0 0
2
43001.6 20
0
14 Logic Display~
6 1552 1300 0 1 2
10 51
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L33
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7743 0 0
2
43001.6 21
0
14 Logic Display~
6 1552 1325 0 1 2
10 15
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L32
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9840 0 0
2
43001.6 22
0
14 Logic Display~
6 1552 1351 0 1 2
10 14
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L31
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6910 0 0
2
43001.6 23
0
14 Logic Display~
6 1552 1274 0 1 2
10 57
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L30
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
449 0 0
2
43001.6 24
0
7 74LS164
127 716 1324 0 12 25
0 63 63 4 62 109 110 111 112 57
51 15 14
0
0 0 4848 0
6 74F164
-21 -51 21 -43
3 U20
-14 4 7 12
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
8761 0 0
2
43001.6 25
0
14 Logic Display~
6 1550 1405 0 1 2
10 58
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L21
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
5.89815e-315 5.44487e-315
0
14 Logic Display~
6 1550 1482 0 1 2
10 55
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L23
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7393 0 0
2
5.89815e-315 5.44746e-315
0
14 Logic Display~
6 1550 1456 0 1 2
10 49
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L24
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7699 0 0
2
5.89815e-315 5.45005e-315
0
14 Logic Display~
6 1549 1558 0 1 2
10 59
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L25
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6638 0 0
2
5.89815e-315 5.45264e-315
0
14 Logic Display~
6 1550 1584 0 1 2
10 61
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L26
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
5.89815e-315 5.45523e-315
0
14 Logic Display~
6 1549 1533 0 1 2
10 53
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L27
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9395 0 0
2
5.89815e-315 5.45782e-315
0
14 Logic Display~
6 1549 1507 0 1 2
10 52
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L28
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3303 0 0
2
5.89815e-315 5.46041e-315
0
14 Logic Display~
6 1550 1608 0 1 2
10 64
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L29
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4498 0 0
2
5.89815e-315 5.463e-315
0
14 Logic Display~
6 1550 1431 0 1 2
10 48
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9728 0 0
2
5.89815e-315 5.46559e-315
0
9 Inverter~
13 662 1610 0 2 22
0 16 64
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3789 0 0
2
5.89815e-315 5.46818e-315
0
9 Inverter~
13 662 1509 0 2 22
0 41 52
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3978 0 0
2
5.89815e-315 5.47077e-315
0
9 Inverter~
13 662 1535 0 2 22
0 40 53
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3494 0 0
2
5.89815e-315 5.47207e-315
0
9 Inverter~
13 662 1586 0 2 22
0 38 61
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3507 0 0
2
5.89815e-315 5.47336e-315
0
9 Inverter~
13 662 1560 0 2 22
0 39 59
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
5151 0 0
2
5.89815e-315 5.47466e-315
0
9 Inverter~
13 663 1458 0 2 22
0 43 49
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3701 0 0
2
5.89815e-315 5.47595e-315
0
9 Inverter~
13 663 1484 0 2 22
0 42 55
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8585 0 0
2
5.89815e-315 5.47725e-315
0
9 Inverter~
13 663 1433 0 2 22
0 44 48
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
8809 0 0
2
5.89815e-315 5.47854e-315
0
9 Inverter~
13 663 1407 0 2 22
0 45 58
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
5993 0 0
2
5.89815e-315 5.47984e-315
0
7 74LS154
95 551 1316 0 22 45
0 2 2 34 35 36 37 113 114 115
116 117 118 16 38 39 40 41 42 43
44 45 119
0
0 0 4848 270
6 74F154
-21 -87 21 -79
3 U17
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
8654 0 0
2
5.89815e-315 5.48113e-315
0
9 4-In NOR~
219 1422 275 0 5 22
0 68 67 66 65 19
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 1 0
1 U
7223 0 0
2
5.89815e-315 5.48243e-315
0
7 74LS126
116 1089 430 0 12 25
0 6 69 6 70 6 71 6 72 27
26 25 24
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
3 U15
-10 -52 11 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3641 0 0
2
5.89815e-315 5.48372e-315
0
7 Ground~
168 1108 510 0 1 3
0 2
0
0 0 53360 270
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3104 0 0
2
5.89815e-315 5.48502e-315
0
7 74LS181
132 1190 471 0 22 45
0 73 49 74 73 65 66 67 68 78
77 76 75 48 2 120 121 122 123 69
70 71 72
0
0 0 4848 180
7 74LS181
-24 -69 25 -61
3 U14
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
3296 0 0
2
5.89815e-315 5.48631e-315
0
6 PROM32
80 777 600 0 14 29
0 10 2 23 22 21 20 31 30 29
28 27 26 25 24
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8534 0 0
2
5.89815e-315 5.48761e-315
0
BKGAJAEAFAGAHIILJAAAAFCAAAAAAAAFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 Ground~
168 389 599 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
949 0 0
2
5.89815e-315 5.4889e-315
0
7 74LS173
129 771 440 0 14 29
0 2 11 11 3 24 25 26 27 2
2 79 80 81 82
0
0 0 4848 270
6 74F173
-21 -51 21 -43
3 U12
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3371 0 0
2
5.89815e-315 5.4902e-315
0
7 Ground~
168 869 405 0 1 3
0 2
0
0 0 53360 90
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7311 0 0
2
5.89815e-315 5.49149e-315
0
7 Ground~
168 546 479 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
5.89815e-315 5.49279e-315
0
7 74LS257
147 614 517 0 14 29
0 83 79 84 80 85 81 86 82 87
2 20 21 22 23
0
0 0 4848 270
6 74F257
-21 -60 21 -52
3 U11
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3526 0 0
2
5.89815e-315 5.49408e-315
0
7 Ground~
168 475 168 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4129 0 0
2
5.89815e-315 5.49538e-315
0
2 +V
167 598 114 0 1 3
0 88
0
0 0 54256 0
2 5V
-8 -22 6 -14
3 V17
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6278 0 0
2
5.89815e-315 5.49667e-315
0
7 74LS193
137 663 168 0 14 29
0 15 88 12 2 27 26 25 24 124
125 92 91 90 89
0
0 0 4848 0
6 74F193
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3482 0 0
2
5.89815e-315 5.49797e-315
0
7 74LS126
116 826 169 0 12 25
0 14 92 14 91 14 90 14 89 27
26 25 24
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
8323 0 0
2
5.89815e-315 5.49926e-315
0
7 74LS126
116 845 1176 0 12 25
0 13 97 13 98 13 99 13 100 24
25 26 27
0
0 0 4848 0
6 74F126
-21 -51 21 -43
2 U8
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3984 0 0
2
5.89815e-315 5.50056e-315
0
7 Ground~
168 743 1174 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7622 0 0
2
5.89815e-315 5.50185e-315
0
7 74LS173
129 671 1128 0 14 29
0 2 18 18 3 24 25 26 27 2
2 97 98 99 100
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U7
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
816 0 0
2
5.89815e-315 5.50315e-315
0
7 74LS173
129 542 1127 0 14 29
0 17 18 18 3 28 29 30 31 2
2 37 36 35 34
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U6
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4656 0 0
2
5.89815e-315 5.50444e-315
0
14 Logic Display~
6 1390 1160 0 1 2
10 104
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6356 0 0
2
5.89815e-315 5.50574e-315
0
14 Logic Display~
6 1370 1160 0 1 2
10 103
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7479 0 0
2
5.89815e-315 5.50703e-315
0
14 Logic Display~
6 1350 1160 0 1 2
10 102
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5690 0 0
2
5.89815e-315 5.50833e-315
0
14 Logic Display~
6 1331 1160 0 1 2
10 101
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5617 0 0
2
5.89815e-315 5.50963e-315
0
7 Ground~
168 1253 1131 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3903 0 0
2
5.89815e-315 5.51092e-315
0
7 74LS173
129 1158 1090 0 14 29
0 2 5 5 3 27 26 25 24 2
2 101 102 103 104
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U5
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4452 0 0
2
5.89815e-315 5.51222e-315
0
7 Ground~
168 1400 746 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6282 0 0
2
5.89815e-315 5.51286e-315
0
7 74LS126
116 1090 852 0 12 25
0 7 93 7 94 7 95 7 96 27
26 25 24
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
7187 0 0
2
5.89815e-315 5.51351e-315
0
7 74LS257
147 1323 708 0 14 29
0 33 93 108 94 107 95 106 96 105
2 78 77 76 75
0
0 0 4848 90
6 74F257
-21 -60 21 -52
2 U3
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
6866 0 0
2
5.89815e-315 5.51416e-315
0
7 74LS126
116 1091 294 0 12 25
0 9 65 9 66 9 67 9 68 27
26 25 24
0
0 0 4848 180
7 74LS126
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
7670 0 0
2
5.89815e-315 5.51481e-315
0
7 Ground~
168 1254 242 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
951 0 0
2
5.89815e-315 5.51545e-315
0
7 74LS173
129 1159 200 0 14 29
0 2 8 8 3 27 26 25 24 2
2 65 66 67 68
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U1
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
9536 0 0
2
5.89815e-315 5.5161e-315
0
14 Logic Display~
6 916 1239 0 1 2
10 31
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L16
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5495 0 0
2
43001.6 26
0
14 Logic Display~
6 935 1239 0 1 2
10 30
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L15
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8152 0 0
2
43001.6 27
0
14 Logic Display~
6 955 1239 0 1 2
10 29
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L14
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6223 0 0
2
43001.6 28
0
14 Logic Display~
6 975 1239 0 1 2
10 28
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L13
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5441 0 0
2
43001.6 29
0
14 Logic Display~
6 1053 1239 0 1 2
10 24
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L12
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3189 0 0
2
43001.6 30
0
14 Logic Display~
6 1033 1239 0 1 2
10 25
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L11
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8460 0 0
2
43001.6 31
0
14 Logic Display~
6 1013 1239 0 1 2
10 26
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L10
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5179 0 0
2
43001.6 32
0
14 Logic Display~
6 994 1239 0 1 2
10 27
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
43001.6 33
0
14 Logic Display~
6 994 94 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3928 0 0
2
43001.6 34
0
14 Logic Display~
6 1013 94 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
363 0 0
2
43001.6 35
0
14 Logic Display~
6 1033 94 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8132 0 0
2
43001.6 36
0
14 Logic Display~
6 1053 94 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
65 0 0
2
43001.6 37
0
14 Logic Display~
6 975 94 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6609 0 0
2
43001.6 38
0
14 Logic Display~
6 955 94 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8995 0 0
2
43001.6 39
0
14 Logic Display~
6 935 94 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3918 0 0
2
43001.6 40
0
14 Logic Display~
6 916 94 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7519 0 0
2
43001.6 41
0
273
2 0 3 0 0 4096 0 27 0 0 17 2
313 1209
169 1209
3 3 4 0 0 8320 0 27 57 0 0 5
358 1200
358 1227
660 1227
660 1324
684 1324
1 0 5 0 0 8320 0 17 0 0 59 5
1281 1947
1799 1947
1799 1111
1534 1111
1534 1031
1 0 6 0 0 8192 0 18 0 0 124 4
1156 1950
1156 1927
1630 1927
1630 1829
1 0 7 0 0 8192 0 19 0 0 188 4
1024 1947
1024 1916
1560 1916
1560 1835
1 0 8 0 0 8192 0 20 0 0 257 4
899 1945
899 1894
1136 1894
1136 1840
1 0 9 0 0 8192 0 21 0 0 247 4
776 1953
776 1866
1414 1866
1414 1712
1 0 10 0 0 4096 0 22 0 0 26 4
660 1960
660 1833
771 1833
771 1799
1 0 11 0 0 4096 0 23 0 0 62 2
560 1962
560 1781
1 0 12 0 0 4096 0 24 0 0 171 2
473 1960
473 1775
1 0 13 0 0 4096 0 25 0 0 196 2
384 1963
384 1794
1 0 14 0 0 4096 0 26 0 0 180 2
289 1963
289 1632
1 0 15 0 0 4096 0 16 0 0 87 2
174 1962
174 1637
1 0 15 0 0 4096 0 15 0 0 206 2
74 1969
74 1625
1 0 16 0 0 4096 0 27 0 0 16 2
313 1191
267 1191
0 0 16 0 0 8320 0 0 0 47 0 3
562 1599
267 1599
267 1176
0 0 3 0 0 8192 0 0 0 218 64 3
167 1020
169 1020
169 1230
2 0 14 0 0 4096 0 28 0 0 101 3
398 1388
776 1388
776 1355
3 1 17 0 0 8320 0 28 94 0 0 5
389 1339
389 1201
610 1201
610 1097
571 1097
1 1 2 0 0 4096 0 28 29 0 0 2
380 1388
380 1386
9 0 2 0 0 4096 0 94 0 0 213 2
571 1167
571 1175
0 0 18 0 0 4096 0 0 0 41 205 3
554 1065
469 1065
469 1075
1 0 2 0 0 0 0 30 0 0 112 2
571 1271
571 1272
1 5 19 0 0 12416 0 50 77 0 0 5
791 1639
791 1260
1486 1260
1486 275
1461 275
6 11 20 0 0 4224 0 81 86 0 0 3
745 636
631 636
631 554
3 1 10 0 0 20608 0 31 81 0 0 9
937 1790
937 1799
710 1799
710 1374
785 1374
785 650
731 650
731 564
739 564
5 12 21 0 0 4224 0 81 86 0 0 3
745 627
613 627
613 554
13 4 22 0 0 8320 0 86 81 0 0 3
595 554
595 618
745 618
14 3 23 0 0 8320 0 86 81 0 0 3
577 554
577 609
745 609
0 14 24 0 0 4096 0 0 81 266 0 2
1053 636
809 636
0 13 25 0 0 4096 0 0 81 267 0 2
1033 627
809 627
0 12 26 0 0 4096 0 0 81 268 0 2
1013 618
809 618
0 11 27 0 0 4096 0 0 81 269 0 2
994 609
809 609
0 10 28 0 0 4096 0 0 81 270 0 2
975 600
809 600
0 9 29 0 0 4096 0 0 81 271 0 2
955 591
809 591
0 8 30 0 0 4096 0 0 81 272 0 2
935 582
809 582
0 7 31 0 0 4096 0 0 81 273 0 2
916 573
809 573
1 2 2 0 0 4224 0 82 81 0 0 2
396 600
745 600
0 2 12 0 0 4096 0 0 31 171 0 4
614 1775
893 1775
893 1745
928 1745
1 3 32 0 0 4224 0 31 33 0 0 3
946 1745
946 1747
945 1747
3 2 18 0 0 0 0 94 94 0 0 5
553 1091
554 1091
554 1065
562 1065
562 1091
2 1 33 0 0 4224 0 32 103 0 0 3
1761 762
1282 762
1282 739
14 3 34 0 0 4224 0 94 76 0 0 4
508 1161
508 1257
535 1257
535 1286
13 4 35 0 0 4224 0 94 76 0 0 4
517 1161
517 1262
526 1262
526 1286
12 5 36 0 0 4224 0 94 76 0 0 4
526 1161
526 1267
517 1267
517 1286
11 6 37 0 0 4224 0 94 76 0 0 4
535 1161
535 1272
508 1272
508 1286
13 1 16 0 0 0 0 76 67 0 0 3
562 1356
562 1610
647 1610
14 1 38 0 0 4224 0 76 70 0 0 3
553 1356
553 1586
647 1586
15 1 39 0 0 4224 0 76 71 0 0 3
544 1356
544 1560
647 1560
16 1 40 0 0 4224 0 76 69 0 0 3
535 1356
535 1535
647 1535
17 1 41 0 0 4224 0 76 68 0 0 3
526 1356
526 1509
647 1509
18 1 42 0 0 8320 0 76 73 0 0 3
517 1356
517 1484
648 1484
19 1 43 0 0 8320 0 76 72 0 0 3
508 1356
508 1458
648 1458
20 1 44 0 0 8320 0 76 74 0 0 3
499 1356
499 1433
648 1433
21 1 45 0 0 8320 0 76 75 0 0 3
490 1356
490 1407
648 1407
2 3 46 0 0 4224 0 35 47 0 0 3
987 1799
987 1689
955 1689
3 1 46 0 0 0 0 47 33 0 0 4
955 1689
955 1694
954 1694
954 1695
1 0 2 0 0 0 0 100 0 0 224 3
1187 1060
1225 1060
1225 1132
2 3 5 0 0 128 0 34 100 0 0 3
1684 1031
1169 1031
1169 1054
0 1 9 0 0 0 0 0 34 247 0 3
1950 1033
1720 1033
1720 1031
1 0 13 0 0 0 0 37 0 0 196 4
866 1700
866 1699
875 1699
875 1685
3 2 11 0 0 12416 0 37 83 0 0 6
857 1752
857 1781
14 1781
14 295
791 295
791 404
3 2 47 0 0 4224 0 49 38 0 0 3
773 1732
773 1743
764 1743
0 1 3 0 0 0 0 0 2 0 0 3
167 1225
169 1225
169 1396
1 0 48 0 0 4096 0 39 0 0 134 2
1875 587
1875 634
0 1 49 0 0 4096 0 0 40 243 0 3
1934 764
1934 545
1873 545
4 2 50 0 0 8320 0 45 41 0 0 3
1032 1670
1084 1670
1084 1765
1 0 51 0 0 4096 0 41 0 0 99 2
1102 1765
1102 1304
1 0 52 0 0 4096 0 42 0 0 106 2
1192 1722
1192 1511
2 0 51 0 0 0 0 42 0 0 99 2
1174 1722
1174 1304
1 0 51 0 0 0 0 43 0 0 99 2
1134 1667
1134 1304
2 0 53 0 0 4096 0 43 0 0 105 2
1116 1667
1116 1537
1 0 52 0 0 0 0 44 0 0 106 2
1051 1680
1051 1511
3 1 54 0 0 4224 0 44 46 0 0 4
1042 1726
1042 1742
1033 1742
1033 1743
2 4 50 0 0 0 0 44 45 0 0 3
1033 1680
1033 1670
1032 1670
1 0 55 0 0 4096 0 45 0 0 107 2
1041 1624
1041 1486
2 0 49 0 0 0 0 45 0 0 108 2
1032 1625
1032 1460
3 0 48 0 0 4096 0 45 0 0 109 2
1023 1624
1023 1435
2 0 51 0 0 0 0 46 0 0 99 2
1015 1743
1015 1304
3 1 56 0 0 8320 0 46 35 0 0 4
1024 1788
1024 1796
1005 1796
1005 1799
2 0 15 0 0 4096 0 33 0 0 100 4
936 1695
936 1344
937 1344
937 1329
2 0 57 0 0 4096 0 47 0 0 98 2
946 1644
946 1278
1 0 58 0 0 4096 0 47 0 0 110 2
964 1644
964 1409
2 0 14 0 0 0 0 37 0 0 101 4
848 1700
848 1370
857 1370
857 1355
1 0 51 0 0 0 0 48 0 0 99 2
884 1640
884 1304
2 0 58 0 0 0 0 48 0 0 110 2
866 1640
866 1409
0 1 15 0 0 12416 0 0 89 100 0 7
825 1329
825 1637
6 1637
6 110
385 110
385 141
631 141
1 0 51 0 0 0 0 38 0 0 99 5
764 1761
791 1761
791 1730
820 1730
820 1304
2 0 59 0 0 4096 0 49 0 0 104 2
764 1686
764 1562
1 3 60 0 0 4224 0 49 50 0 0 2
782 1686
782 1684
2 0 61 0 0 4096 0 50 0 0 103 2
773 1639
773 1588
1 4 62 0 0 8320 0 51 57 0 0 3
675 1357
678 1357
678 1342
3 0 51 0 0 0 0 52 0 0 99 3
736 1252
779 1252
779 1304
2 0 15 0 0 0 0 52 0 0 100 3
735 1261
774 1261
774 1329
1 0 14 0 0 0 0 52 0 0 101 3
736 1270
770 1270
770 1355
2 0 63 0 0 4096 0 57 0 0 97 3
684 1306
669 1306
669 1297
1 4 63 0 0 8320 0 57 52 0 0 4
684 1297
669 1297
669 1261
684 1261
9 1 57 0 0 12416 0 57 56 0 0 4
748 1333
766 1333
766 1278
1536 1278
10 1 51 0 0 12416 0 57 53 0 0 4
748 1342
759 1342
759 1304
1536 1304
1 11 15 0 0 0 0 54 57 0 0 4
1536 1329
754 1329
754 1351
748 1351
1 12 14 0 0 4096 0 55 57 0 0 4
1536 1355
754 1355
754 1360
748 1360
2 1 64 0 0 8320 0 67 65 0 0 3
683 1610
683 1612
1534 1612
2 1 61 0 0 8320 0 70 62 0 0 3
683 1586
683 1588
1534 1588
2 1 59 0 0 8320 0 71 61 0 0 3
683 1560
683 1562
1533 1562
2 1 53 0 0 8320 0 69 63 0 0 3
683 1535
683 1537
1533 1537
2 1 52 0 0 8320 0 68 64 0 0 3
683 1509
683 1511
1533 1511
2 1 55 0 0 8320 0 73 59 0 0 3
684 1484
684 1486
1534 1486
2 1 49 0 0 8192 0 72 60 0 0 3
684 1458
684 1460
1534 1460
2 1 48 0 0 8192 0 74 66 0 0 3
684 1433
684 1435
1534 1435
2 1 58 0 0 8320 0 75 58 0 0 3
684 1407
684 1409
1534 1409
0 2 64 0 0 0 0 0 67 0 0 4
684 1610
682 1610
682 1610
683 1610
1 2 2 0 0 0 0 76 76 0 0 4
571 1280
571 1272
562 1272
562 1280
0 4 65 0 0 4096 0 0 77 120 0 4
1233 316
1356 316
1356 289
1405 289
0 3 66 0 0 4096 0 0 77 119 0 4
1245 299
1343 299
1343 280
1405 280
0 2 67 0 0 4096 0 0 77 118 0 4
1255 282
1334 282
1334 271
1405 271
0 1 68 0 0 4096 0 0 77 117 0 2
1265 262
1405 262
8 8 68 0 0 8320 0 80 104 0 0 4
1228 457
1265 457
1265 262
1123 262
7 0 67 0 0 8320 0 80 0 0 254 4
1228 466
1255 466
1255 280
1134 280
6 0 66 0 0 8320 0 80 0 0 253 4
1228 475
1245 475
1245 298
1143 298
0 5 65 0 0 8320 0 0 80 252 0 4
1152 316
1236 316
1236 484
1228 484
7 0 6 0 0 0 0 78 0 0 124 2
1121 407
1128 407
5 0 6 0 0 0 0 78 0 0 124 2
1121 425
1128 425
3 0 6 0 0 0 0 78 0 0 124 2
1121 443
1128 443
3 1 6 0 0 12416 0 41 78 0 0 7
1093 1810
1093 1829
1939 1829
1939 375
1128 375
1128 461
1121 461
2 19 69 0 0 4224 0 78 80 0 0 3
1121 452
1152 452
1152 448
4 20 70 0 0 4224 0 78 80 0 0 4
1121 434
1147 434
1147 439
1152 439
6 21 71 0 0 4224 0 78 80 0 0 4
1121 416
1142 416
1142 430
1152 430
22 8 72 0 0 12416 0 80 78 0 0 4
1152 421
1146 421
1146 398
1121 398
9 0 27 0 0 0 0 78 0 0 269 2
1057 452
994 452
10 0 26 0 0 0 0 78 0 0 268 2
1057 434
1013 434
11 0 25 0 0 0 0 78 0 0 267 2
1057 416
1033 416
12 0 24 0 0 0 0 78 0 0 266 2
1057 398
1053 398
14 1 2 0 0 0 0 80 79 0 0 2
1158 511
1115 511
13 0 48 0 0 16512 0 80 0 0 109 7
1158 520
1146 520
1146 634
1929 634
1929 1817
1231 1817
1231 1435
4 2 73 0 0 4224 0 80 40 0 0 4
1222 493
1839 493
1839 545
1837 545
3 2 74 0 0 4224 0 80 39 0 0 4
1222 502
1807 502
1807 587
1839 587
2 0 49 0 0 0 0 80 0 0 66 4
1222 511
1776 511
1776 561
1934 561
1 2 73 0 0 0 0 80 40 0 0 4
1222 520
1743 520
1743 545
1837 545
12 14 75 0 0 8320 0 80 103 0 0 3
1228 421
1354 421
1354 675
11 13 76 0 0 8320 0 80 103 0 0 3
1228 430
1336 430
1336 675
10 12 77 0 0 8320 0 80 103 0 0 3
1228 439
1318 439
1318 675
9 11 78 0 0 8320 0 80 103 0 0 3
1228 448
1300 448
1300 675
8 0 31 0 0 8192 0 94 0 0 273 3
508 1097
508 935
916 935
0 7 30 0 0 4096 0 0 94 272 0 3
935 946
517 946
517 1097
6 0 29 0 0 8192 0 94 0 0 271 3
526 1097
526 961
955 961
5 0 28 0 0 8192 0 94 0 0 270 3
535 1097
535 975
975 975
2 11 79 0 0 8320 0 86 83 0 0 4
640 490
640 483
764 483
764 474
12 4 80 0 0 8320 0 83 86 0 0 4
755 474
755 480
622 480
622 490
6 13 81 0 0 8320 0 86 83 0 0 4
604 490
604 477
746 477
746 474
14 8 82 0 0 4224 0 83 86 0 0 3
737 474
586 474
586 490
4 0 3 0 0 8192 0 83 0 0 218 3
773 410
773 275
167 275
5 0 24 0 0 8192 0 83 0 0 266 3
764 410
764 363
1053 363
6 0 25 0 0 8192 0 83 0 0 267 3
755 410
755 353
1033 353
7 0 26 0 0 8192 0 83 0 0 268 3
746 410
746 342
1013 342
8 0 27 0 0 8192 0 83 0 0 269 3
737 410
737 330
994 330
3 0 11 0 0 0 0 83 0 0 62 3
782 404
782 395
791 395
9 0 2 0 0 0 0 83 0 0 158 2
800 480
800 490
10 0 2 0 0 0 0 83 0 0 159 4
791 480
791 490
851 490
851 406
1 1 2 0 0 0 0 83 84 0 0 3
800 410
800 406
862 406
1 10 2 0 0 0 0 85 86 0 0 3
553 480
568 480
568 484
1 1 83 0 0 8320 0 86 1 0 0 5
649 490
649 359
263 359
263 441
218 441
1 3 84 0 0 8320 0 3 86 0 0 4
381 488
381 412
631 412
631 490
1 5 85 0 0 8320 0 4 86 0 0 4
349 487
349 397
613 397
613 490
1 7 86 0 0 8320 0 5 86 0 0 4
318 487
318 383
595 383
595 490
1 9 87 0 0 8320 0 6 86 0 0 4
285 485
285 370
577 370
577 490
9 0 27 0 0 0 0 90 0 0 269 2
858 151
994 151
10 0 26 0 0 0 0 90 0 0 268 2
858 169
1013 169
11 0 25 0 0 0 0 90 0 0 267 2
858 187
1033 187
12 0 24 0 0 0 0 90 0 0 266 2
858 205
1053 205
1 4 2 0 0 0 0 87 89 0 0 3
482 169
482 168
631 168
3 3 12 0 0 12416 0 89 38 0 0 7
625 159
625 158
2 158
2 1775
616 1775
616 1752
713 1752
2 1 88 0 0 4224 0 89 88 0 0 3
631 150
598 150
598 123
0 5 27 0 0 4096 0 0 89 269 0 4
994 248
593 248
593 177
631 177
0 6 26 0 0 4096 0 0 89 268 0 4
1013 240
602 240
602 186
631 186
0 7 25 0 0 4096 0 0 89 267 0 4
1033 231
611 231
611 195
631 195
0 8 24 0 0 4096 0 0 89 266 0 4
1053 222
620 222
620 204
631 204
1 0 14 0 0 0 0 90 0 0 180 2
794 142
780 142
3 0 14 0 0 0 0 90 0 0 180 2
794 160
780 160
5 0 14 0 0 0 0 90 0 0 180 2
794 178
780 178
0 7 14 0 0 12416 0 0 90 101 0 7
830 1355
830 1632
10 1632
10 68
780 68
780 196
794 196
8 14 89 0 0 8320 0 90 89 0 0 3
794 205
794 204
695 204
6 13 90 0 0 12416 0 90 89 0 0 4
794 187
748 187
748 195
695 195
4 12 91 0 0 4224 0 90 89 0 0 4
794 169
740 169
740 186
695 186
11 2 92 0 0 12416 0 89 90 0 0 4
695 177
731 177
731 151
794 151
7 0 7 0 0 0 0 102 0 0 188 2
1122 829
1148 829
5 0 7 0 0 0 0 102 0 0 188 2
1122 847
1148 847
3 0 7 0 0 0 0 102 0 0 188 2
1122 865
1148 865
3 1 7 0 0 12416 0 42 102 0 0 7
1183 1767
1183 1835
1945 1835
1945 802
1148 802
1148 883
1122 883
2 0 93 0 0 4096 0 102 0 0 242 2
1122 874
1290 874
4 0 94 0 0 4096 0 102 0 0 241 2
1122 856
1309 856
6 0 95 0 0 4224 0 102 0 0 240 2
1122 838
1327 838
8 0 96 0 0 4224 0 102 0 0 239 2
1122 820
1345 820
7 0 13 0 0 0 0 91 0 0 196 2
813 1203
758 1203
5 0 13 0 0 0 0 91 0 0 196 3
813 1185
813 1171
758 1171
3 0 13 0 0 0 0 91 0 0 196 2
813 1167
758 1167
3 1 13 0 0 12416 0 48 91 0 0 8
875 1685
886 1685
886 1794
26 1794
26 1238
758 1238
758 1149
813 1149
11 2 97 0 0 8320 0 93 91 0 0 5
664 1162
664 1186
793 1186
793 1158
813 1158
12 0 27 0 0 0 0 91 0 0 269 2
877 1212
994 1212
11 0 26 0 0 0 0 91 0 0 268 2
877 1194
1013 1194
10 0 25 0 0 0 0 91 0 0 267 2
877 1176
1033 1176
9 0 24 0 0 0 0 91 0 0 266 2
877 1158
1053 1158
12 4 98 0 0 8320 0 93 91 0 0 5
655 1162
655 1190
807 1190
807 1176
813 1176
13 6 99 0 0 8320 0 93 91 0 0 3
646 1162
646 1194
813 1194
14 8 100 0 0 8320 0 93 91 0 0 3
637 1162
637 1212
813 1212
3 2 18 0 0 8320 0 93 36 0 0 5
682 1092
682 1075
346 1075
346 1059
341 1059
0 1 15 0 0 0 0 0 36 100 0 5
837 1329
837 1625
22 1625
22 1059
305 1059
3 2 18 0 0 0 0 93 93 0 0 2
682 1092
691 1092
0 0 3 0 0 0 0 0 0 209 218 2
673 1087
673 1020
4 4 3 0 0 0 0 93 94 0 0 4
673 1098
673 1085
544 1085
544 1097
1 0 2 0 0 0 0 92 0 0 211 4
736 1175
737 1175
737 1175
736 1175
1 0 2 0 0 0 0 93 0 0 212 4
700 1098
736 1098
736 1175
699 1175
0 9 2 0 0 0 0 0 93 213 0 3
690 1175
700 1175
700 1168
10 10 2 0 0 0 0 94 93 0 0 4
562 1167
562 1175
691 1175
691 1168
5 0 24 0 0 0 0 93 0 0 266 3
664 1098
664 1068
1053 1068
6 0 25 0 0 0 0 93 0 0 267 3
655 1098
655 1063
1033 1063
7 0 26 0 0 0 0 93 0 0 268 3
646 1098
646 1057
1013 1057
8 0 27 0 0 0 0 93 0 0 269 3
637 1098
637 1051
994 1051
4 0 3 0 0 8192 0 100 0 0 261 4
1160 1060
1160 1020
167 1020
167 31
11 1 101 0 0 8320 0 100 98 0 0 4
1151 1124
1151 1217
1331 1217
1331 1178
12 1 102 0 0 8320 0 100 97 0 0 4
1142 1124
1142 1210
1350 1210
1350 1178
13 1 103 0 0 8320 0 100 96 0 0 4
1133 1124
1133 1199
1370 1199
1370 1178
14 1 104 0 0 8320 0 100 95 0 0 4
1124 1124
1124 1189
1390 1189
1390 1178
9 0 2 0 0 0 0 100 0 0 224 2
1187 1130
1187 1132
10 1 2 0 0 0 0 100 99 0 0 3
1178 1130
1178 1132
1246 1132
2 0 5 0 0 0 0 100 0 0 59 2
1178 1054
1178 1031
5 0 27 0 0 0 0 100 0 0 269 3
1151 1060
1151 1036
994 1036
6 0 26 0 0 0 0 100 0 0 268 3
1142 1060
1142 1042
1013 1042
7 0 25 0 0 0 0 100 0 0 267 3
1133 1060
1133 1050
1033 1050
8 0 24 0 0 0 0 100 0 0 266 2
1124 1060
1053 1060
1 10 2 0 0 0 0 101 103 0 0 3
1393 747
1393 745
1363 745
9 0 27 0 0 0 0 102 0 0 269 2
1058 874
994 874
10 0 26 0 0 0 0 102 0 0 268 2
1058 856
1013 856
11 0 25 0 0 0 0 102 0 0 267 2
1058 838
1033 838
12 0 24 0 0 0 0 102 0 0 266 2
1058 820
1053 820
9 1 105 0 0 8320 0 103 10 0 0 4
1354 739
1354 835
1633 835
1633 955
7 1 106 0 0 8320 0 103 9 0 0 4
1336 739
1336 849
1601 849
1601 954
5 1 107 0 0 8320 0 103 8 0 0 4
1318 739
1318 864
1570 864
1570 954
3 1 108 0 0 8320 0 103 7 0 0 4
1300 739
1300 878
1537 878
1537 952
8 1 96 0 0 0 0 103 11 0 0 4
1345 739
1345 918
1386 918
1386 953
6 1 95 0 0 0 0 103 12 0 0 4
1327 739
1327 928
1354 928
1354 952
4 1 94 0 0 4224 0 103 13 0 0 4
1309 739
1309 938
1323 938
1323 952
2 1 93 0 0 8320 0 103 14 0 0 3
1291 739
1290 739
1290 950
0 1 49 0 0 12416 0 0 32 108 0 5
1222 1460
1222 1824
1934 1824
1934 762
1797 762
0 7 9 0 0 0 0 0 104 245 0 3
1129 290
1129 271
1123 271
0 5 9 0 0 0 0 0 104 246 0 3
1129 307
1129 289
1123 289
3 0 9 0 0 0 0 104 0 0 247 3
1123 307
1129 307
1129 325
1 3 9 0 0 8320 0 104 43 0 0 4
1123 325
1950 325
1950 1712
1125 1712
9 0 27 0 0 0 0 104 0 0 269 2
1059 316
994 316
10 0 26 0 0 0 0 104 0 0 268 2
1059 298
1013 298
11 0 25 0 0 0 0 104 0 0 267 2
1059 280
1033 280
12 0 24 0 0 0 0 104 0 0 266 2
1059 262
1053 262
11 2 65 0 0 0 0 106 104 0 0 3
1152 234
1152 316
1123 316
12 4 66 0 0 0 0 106 104 0 0 3
1143 234
1143 298
1123 298
13 6 67 0 0 0 0 106 104 0 0 3
1134 234
1134 280
1123 280
14 8 68 0 0 0 0 106 104 0 0 3
1125 234
1123 234
1123 262
2 0 8 0 0 0 0 106 0 0 257 2
1179 164
1179 141
3 3 8 0 0 16512 0 35 106 0 0 7
996 1851
1016 1851
1016 1840
1955 1840
1955 141
1170 141
1170 164
1 0 2 0 0 0 0 106 0 0 260 3
1188 170
1220 170
1220 243
9 0 2 0 0 0 0 106 0 0 260 2
1188 240
1188 243
10 1 2 0 0 0 0 106 105 0 0 3
1179 240
1179 243
1247 243
0 4 3 0 0 4224 0 0 106 0 0 3
112 31
1161 31
1161 170
5 0 27 0 0 0 0 106 0 0 269 3
1152 170
1152 146
994 146
6 0 26 0 0 0 0 106 0 0 268 3
1143 170
1143 152
1013 152
7 0 25 0 0 0 0 106 0 0 267 3
1134 170
1134 160
1033 160
8 0 24 0 0 0 0 106 0 0 266 2
1125 170
1053 170
1 1 24 0 0 4224 0 118 111 0 0 2
1053 112
1053 1225
1 1 25 0 0 4224 0 117 112 0 0 2
1033 112
1033 1225
1 1 26 0 0 4224 0 116 113 0 0 2
1013 112
1013 1225
1 1 27 0 0 4224 0 115 114 0 0 2
994 112
994 1225
1 1 28 0 0 4224 0 119 110 0 0 2
975 112
975 1225
1 1 29 0 0 4224 0 120 109 0 0 2
955 112
955 1225
1 1 30 0 0 4224 0 121 108 0 0 2
935 112
935 1225
1 1 31 0 0 4224 0 122 107 0 0 2
916 112
916 1225
58
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1256 1971 1299 1986
1270 1983 1284 1994
2 Lo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1129 1974 1172 1989
1143 1986 1157 1997
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
976 1976 1019 1991
990 1987 1004 1998
2 Eb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
867 1971 910 1986
881 1983 895 1994
2 La
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
749 1976 792 1991
763 1987 777 1998
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
633 1989 676 2004
647 2000 661 2011
2 Ce
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
41 2000 86 2015
56 2011 70 2022
2 Li
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
534 1987 579 2002
549 1999 563 2010
2 Lm
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
439 1989 482 2004
453 2000 467 2011
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
359 1991 402 2006
373 2003 387 2014
2 Ei
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
250 1993 293 2008
264 2004 278 2015
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
134 1994 179 2009
149 2006 163 2017
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
190 446 288 469
202 456 275 471
9 SM(MAR=1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
704 1588 755 1611
717 1598 741 1613
3 HLT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
708 1565 751 1588
721 1575 737 1590
2 JZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1537 757 1560
720 1547 744 1562
3 JMP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1514 757 1537
720 1524 744 1539
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
707 1488 758 1511
720 1498 744 1513
3 MOV
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1460 757 1483
720 1470 744 1485
3 AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
706 1436 757 1459
719 1446 743 1461
3 SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1409 757 1432
720 1419 744 1434
3 ADD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
709 1382 758 1405
721 1392 745 1407
3 LDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 1331 833 1354
803 1341 819 1356
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 1304 829 1327
800 1314 816 1329
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
789 1280 832 1303
802 1290 818 1305
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 1252 833 1275
803 1262 819 1277
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1627 119 1664 143
1638 128 1652 144
2 LA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1653 303 1680 327
1658 307 1674 323
2 EA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1661 739 1694 760
1669 746 1685 761
2 RS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1662 778 1695 799
1670 785 1686 800
2 EB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1653 1027 1690 1051
1663 1035 1679 1051
2 LO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
123 41 160 65
133 49 149 65
2 EP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
121 125 158 149
131 133 147 149
2 LP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
119 533 154 555
128 540 144 556
2 CE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
708 78 743 100
717 85 733 101
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
809 364 852 386
818 371 842 387
3 MAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
420 418 527 440
429 425 517 441
11 INPUT & MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
755 652 798 674
764 660 788 676
3 RAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
654 986 689 1008
663 994 679 1010
2 IR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
125 274 162 296
135 281 151 297
2 LM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
130 1058 165 1080
139 1065 155 1081
2 LI
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 1237 168 1259
142 1245 158 1261
2 EI
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
117 7 176 29
126 15 166 31
5 CLOCK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
122 86 157 108
131 93 147 109
2 CP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1647 633 1690 655
1656 640 1680 656
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1750 518 1785 540
1759 525 1775 541
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1782 515 1817 537
1791 523 1807 539
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1813 505 1848 527
1822 512 1838 528
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1714 521 1749 543
1723 529 1739 545
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1645 349 1682 371
1655 356 1671 372
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1275 201 1304 223
1285 208 1293 224
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1373 426 1416 448
1382 434 1406 450
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1409 699 1452 721
1418 706 1442 722
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1163 919 1190 941
1172 926 1180 942
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1504 913 1531 935
1513 920 1521 936
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1229 1051 1304 1073
1238 1058 1294 1074
7 OUT REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1418 1148 1493 1170
1427 1155 1483 1171
7 DISPLAY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
200 1395 265 1418
212 1405 252 1420
5 CLOCK
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
