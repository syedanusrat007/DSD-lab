CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 34 246 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 37 203 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 36 159 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89773e-315 0
0
13 Logic Switch~
5 39 106 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89773e-315 0
0
7 74LS173
129 408 78 0 14 29
0 10 11 12 13 14 15 16 17 18
19 2 3 4 5
0
0 0 4832 0
7 74LS173
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
8157 0 0
2
5.89773e-315 0
0
7 74LS157
122 251 144 0 14 29
0 20 9 5 8 4 7 3 6 2
21 22 23 24 25
0
0 0 4832 0
7 74LS157
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
5572 0 0
2
5.89773e-315 0
0
8
9 11 2 0 0 12416 0 6 5 0 0 6
219 180
189 180
189 16
469 16
469 87
440 87
7 12 3 0 0 12416 0 6 5 0 0 6
219 162
194 162
194 21
464 21
464 96
440 96
5 13 4 0 0 12416 0 6 5 0 0 6
219 144
199 144
199 26
459 26
459 105
440 105
3 14 5 0 0 12416 0 6 5 0 0 6
219 126
209 126
209 31
454 31
454 114
440 114
1 8 6 0 0 4224 0 1 6 0 0 4
46 246
205 246
205 171
219 171
1 6 7 0 0 4224 0 2 6 0 0 4
49 203
200 203
200 153
219 153
1 4 8 0 0 4224 0 3 6 0 0 4
48 159
205 159
205 135
219 135
1 2 9 0 0 4224 0 4 6 0 0 4
51 106
205 106
205 117
219 117
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
205 215 282 239
215 223 271 239
7 2:1 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
354 132 447 156
364 140 436 156
9 Input MAR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
