CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
650 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
77
13 Logic Switch~
5 508 53 0 1 11
0 66
0
0 0 21360 782
2 0V
-6 -21 8 -13
3 V12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3756 0 0
2
42939.8 0
0
13 Logic Switch~
5 465 52 0 1 11
0 45
0
0 0 21360 782
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6760 0 0
2
42939.8 0
0
13 Logic Switch~
5 425 52 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
351 0 0
2
42939.8 0
0
13 Logic Switch~
5 381 54 0 1 11
0 14
0
0 0 21360 782
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5352 0 0
2
42939.8 0
0
13 Logic Switch~
5 336 53 0 10 11
0 67 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
485 0 0
2
42939.8 0
0
13 Logic Switch~
5 296 54 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
452 0 0
2
42939.8 0
0
13 Logic Switch~
5 252 56 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
643 0 0
2
42939.8 0
0
13 Logic Switch~
5 214 53 0 1 11
0 15
0
0 0 21360 782
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5563 0 0
2
42939.8 0
0
13 Logic Switch~
5 170 55 0 10 11
0 62 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
934 0 0
2
42939.8 0
0
13 Logic Switch~
5 121 55 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3240 0 0
2
42939.8 0
0
13 Logic Switch~
5 76 55 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3233 0 0
2
42939.8 0
0
13 Logic Switch~
5 35 56 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3635 0 0
2
42939.8 0
0
14 Logic Display~
6 1712 47 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3547 0 0
2
42939.8 0
0
14 Logic Display~
6 1652 46 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
483 0 0
2
42939.8 0
0
14 Logic Display~
6 1560 48 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6126 0 0
2
42939.8 0
0
14 Logic Display~
6 1447 50 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7368 0 0
2
42939.8 0
0
9 4-In NOR~
219 1554 97 0 5 22
0 5 8 7 6 2
0
0 0 624 90
4 4002
-14 -24 14 -16
4 U16A
30 -2 58 6
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 16 0
1 U
3925 0 0
2
42939.8 0
0
9 2-In XOR~
219 1444 98 0 3 22
0 4 9 3
0
0 0 624 90
6 74LS86
-21 -24 21 -16
4 U15A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
6187 0 0
2
42939.8 0
0
14 Logic Display~
6 1362 42 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5866 0 0
2
42939.8 0
0
14 Logic Display~
6 1321 43 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6650 0 0
2
42939.8 0
0
14 Logic Display~
6 1261 45 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8814 0 0
2
42939.8 0
0
14 Logic Display~
6 1215 45 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4714 0 0
2
42939.8 0
0
14 Logic Display~
6 1153 45 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9875 0 0
2
42939.8 0
0
8 2-In OR~
219 793 1113 0 3 22
0 26 15 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
8220 0 0
2
42939.8 11
0
9 3-In AND~
219 728 1102 0 4 22
0 27 17 16 26
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U13C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 13 0
1 U
3691 0 0
2
42939.8 10
0
9 2-In XOR~
219 645 1078 0 3 22
0 14 11 27
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
5196 0 0
2
42939.8 9
0
9 2-In AND~
219 653 1158 0 3 22
0 14 13 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
6182 0 0
2
42939.8 8
0
9 2-In AND~
219 652 1203 0 3 22
0 12 11 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
6326 0 0
2
42939.8 7
0
8 2-In OR~
219 715 1178 0 3 22
0 25 24 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
3247 0 0
2
42939.8 6
0
9 2-In AND~
219 653 1247 0 3 22
0 10 9 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
5235 0 0
2
42939.8 5
0
9 2-In XOR~
219 894 1145 0 3 22
0 21 20 23
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9260 0 0
2
42939.8 4
0
9 2-In XOR~
219 1018 1173 0 3 22
0 23 22 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
583 0 0
2
42939.8 3
0
9 2-In AND~
219 982 1276 0 3 22
0 23 22 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3471 0 0
2
42939.8 2
0
8 2-In OR~
219 1041 1292 0 3 22
0 19 18 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
7124 0 0
2
42939.8 1
0
9 3-In AND~
219 977 1319 0 4 22
0 21 10 20 18
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 13 0
1 U
6160 0 0
2
42939.8 0
0
9 3-In AND~
219 964 999 0 4 22
0 35 10 34 32
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 13 0
1 U
4732 0 0
2
42939.8 0
0
8 2-In OR~
219 1028 972 0 3 22
0 33 32 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
8836 0 0
2
42939.8 11
0
9 2-In AND~
219 969 956 0 3 22
0 37 36 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3346 0 0
2
42939.8 9
0
9 2-In XOR~
219 1005 853 0 3 22
0 37 36 8
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
8546 0 0
2
42939.8 8
0
9 2-In XOR~
219 881 825 0 3 22
0 35 34 37
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
8607 0 0
2
42939.8 7
0
9 2-In AND~
219 640 927 0 3 22
0 10 31 36
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
5781 0 0
2
42939.8 6
0
8 2-In OR~
219 702 858 0 3 22
0 39 38 34
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
6991 0 0
2
42939.8 5
0
9 2-In AND~
219 639 883 0 3 22
0 28 11 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
9631 0 0
2
42939.8 4
0
9 2-In AND~
219 640 838 0 3 22
0 29 13 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
8381 0 0
2
42939.8 3
0
9 2-In XOR~
219 632 758 0 3 22
0 29 11 41
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6697 0 0
2
42939.8 2
0
9 3-In AND~
219 715 782 0 4 22
0 41 17 16 40
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 2 0
1 U
3463 0 0
2
42939.8 1
0
8 2-In OR~
219 780 793 0 3 22
0 40 30 35
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
9605 0 0
2
42939.8 0
0
8 2-In OR~
219 736 473 0 3 22
0 54 43 49
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
936 0 0
2
42939.8 11
0
9 3-In AND~
219 671 462 0 4 22
0 55 17 16 54
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 2 0
1 U
9813 0 0
2
42939.8 10
0
9 2-In XOR~
219 588 438 0 3 22
0 45 11 55
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5286 0 0
2
42939.8 9
0
9 2-In AND~
219 596 518 0 3 22
0 45 13 53
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
9179 0 0
2
42939.8 8
0
9 2-In AND~
219 595 563 0 3 22
0 44 11 52
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3718 0 0
2
42939.8 7
0
8 2-In OR~
219 658 538 0 3 22
0 53 52 48
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4375 0 0
2
42939.8 6
0
9 2-In AND~
219 596 607 0 3 22
0 10 42 50
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3616 0 0
2
42939.8 5
0
9 2-In XOR~
219 837 505 0 3 22
0 49 48 51
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7808 0 0
2
42939.8 4
0
9 2-In XOR~
219 961 533 0 3 22
0 51 50 7
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7498 0 0
2
42939.8 3
0
9 2-In AND~
219 925 636 0 3 22
0 51 50 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9736 0 0
2
42939.8 2
0
9 2-In AND~
219 926 679 0 3 22
0 49 48 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9454 0 0
2
42939.8 1
0
8 2-In OR~
219 984 652 0 3 22
0 47 46 31
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4639 0 0
2
42939.8 0
0
8 2-In OR~
219 985 331 0 3 22
0 57 56 42
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3831 0 0
2
42939.8 0
0
9 2-In AND~
219 927 358 0 3 22
0 59 58 56
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3538 0 0
2
42939.8 0
0
9 2-In AND~
219 926 315 0 3 22
0 61 60 57
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5949 0 0
2
42939.8 0
0
9 2-In XOR~
219 962 212 0 3 22
0 61 60 6
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7130 0 0
2
42939.8 0
0
9 2-In XOR~
219 838 184 0 3 22
0 59 58 61
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4115 0 0
2
42939.8 0
0
9 2-In AND~
219 597 286 0 3 22
0 10 62 60
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3197 0 0
2
42939.8 0
0
8 2-In OR~
219 659 217 0 3 22
0 64 63 58
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
813 0 0
2
42939.8 0
0
9 2-In AND~
219 596 242 0 3 22
0 65 11 63
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3396 0 0
2
42939.8 0
0
9 2-In AND~
219 597 197 0 3 22
0 66 13 64
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6348 0 0
2
42939.8 0
0
9 Inverter~
13 521 78 0 2 22
0 66 65
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
583 0 0
2
42939.8 0
0
9 Inverter~
13 479 77 0 2 22
0 45 44
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
922 0 0
2
42939.8 0
0
9 Inverter~
13 439 77 0 2 22
0 29 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
4442 0 0
2
42939.8 0
0
9 Inverter~
13 397 78 0 2 22
0 14 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
5893 0 0
2
42939.8 0
0
9 Inverter~
13 135 73 0 2 22
0 13 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3814 0 0
2
42939.8 0
0
9 Inverter~
13 49 74 0 2 22
0 16 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3637 0 0
2
42939.8 0
0
9 2-In XOR~
219 589 117 0 3 22
0 66 11 69
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6890 0 0
2
42939.8 0
0
9 3-In AND~
219 672 141 0 4 22
0 69 17 16 68
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
3933 0 0
2
42939.8 0
0
8 2-In OR~
219 737 152 0 3 22
0 68 67 59
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3432 0 0
2
42939.8 0
0
145
1 5 2 0 0 4224 0 15 17 0 0 2
1560 66
1560 64
1 3 3 0 0 0 0 16 18 0 0 2
1447 68
1447 68
0 1 4 0 0 4096 0 0 13 11 0 3
1153 259
1712 259
1712 65
0 1 5 0 0 4096 0 0 14 12 0 3
1215 229
1652 229
1652 64
0 4 6 0 0 4096 0 0 17 96 0 3
1362 181
1574 181
1574 120
0 3 7 0 0 4096 0 0 17 14 0 3
1321 168
1565 168
1565 120
0 2 8 0 0 4096 0 0 17 13 0 3
1261 151
1556 151
1556 120
0 1 5 0 0 0 0 0 17 12 0 3
1215 133
1547 133
1547 120
2 0 9 0 0 4224 0 18 0 0 26 3
1456 117
1456 1058
1090 1058
1 0 4 0 0 0 0 18 0 0 11 2
1438 117
1153 117
0 1 4 0 0 4224 0 0 23 27 0 2
1153 1292
1153 63
3 1 5 0 0 8320 0 32 22 0 0 3
1051 1173
1215 1173
1215 63
3 1 8 0 0 8320 0 39 21 0 0 3
1038 853
1261 853
1261 63
3 1 7 0 0 8320 0 56 20 0 0 3
994 533
1321 533
1321 61
2 0 10 0 0 4096 0 35 0 0 127 2
953 1319
70 1319
1 0 10 0 0 0 0 30 0 0 127 2
629 1238
70 1238
2 0 11 0 0 4096 0 28 0 0 144 2
628 1212
76 1212
1 0 12 0 0 4096 0 28 0 0 125 2
628 1194
418 1194
2 0 13 0 0 4096 0 27 0 0 143 2
629 1167
121 1167
1 0 14 0 0 4096 0 27 0 0 137 2
629 1149
381 1149
2 0 15 0 0 4096 0 24 0 0 141 2
780 1122
214 1122
3 0 16 0 0 4096 0 25 0 0 145 2
704 1111
35 1111
2 0 17 0 0 4096 0 25 0 0 126 2
704 1102
156 1102
2 0 11 0 0 4096 0 26 0 0 144 2
629 1087
76 1087
1 0 14 0 0 0 0 26 0 0 137 2
629 1069
381 1069
0 2 9 0 0 0 0 0 30 54 0 5
1090 972
1090 1348
614 1348
614 1256
629 1256
3 0 4 0 0 0 0 34 0 0 0 2
1074 1292
1197 1292
4 2 18 0 0 12416 0 35 34 0 0 4
998 1319
1004 1319
1004 1301
1028 1301
3 1 19 0 0 4224 0 33 34 0 0 4
1003 1276
1021 1276
1021 1283
1028 1283
0 3 20 0 0 8320 0 0 35 36 0 3
797 1178
797 1328
953 1328
0 1 21 0 0 4224 0 0 35 37 0 3
839 1113
839 1310
953 1310
0 2 22 0 0 8192 0 0 33 34 0 3
897 1247
897 1285
958 1285
1 0 23 0 0 8320 0 33 0 0 35 3
958 1267
939 1267
939 1145
3 2 22 0 0 4224 0 30 32 0 0 4
674 1247
986 1247
986 1182
1002 1182
3 1 23 0 0 0 0 31 32 0 0 3
927 1145
1002 1145
1002 1164
3 2 20 0 0 0 0 29 31 0 0 4
748 1178
871 1178
871 1154
878 1154
3 1 21 0 0 0 0 24 31 0 0 4
826 1113
859 1113
859 1136
878 1136
3 2 24 0 0 8320 0 28 29 0 0 3
673 1203
673 1187
702 1187
3 1 25 0 0 8320 0 27 29 0 0 3
674 1158
674 1169
702 1169
4 1 26 0 0 8320 0 25 24 0 0 3
749 1102
749 1104
780 1104
3 1 27 0 0 4224 0 26 25 0 0 4
678 1078
695 1078
695 1093
704 1093
2 0 10 0 0 0 0 36 0 0 127 2
940 999
70 999
1 0 10 0 0 0 0 41 0 0 127 2
616 918
70 918
2 0 11 0 0 0 0 43 0 0 144 2
615 892
76 892
1 0 28 0 0 4096 0 43 0 0 124 2
615 874
460 874
2 0 13 0 0 0 0 44 0 0 143 2
616 847
121 847
1 0 29 0 0 4096 0 44 0 0 136 2
616 829
425 829
2 0 30 0 0 4096 0 47 0 0 140 2
767 802
252 802
3 0 16 0 0 0 0 46 0 0 145 2
691 791
35 791
2 0 17 0 0 0 0 46 0 0 126 2
691 782
156 782
2 0 11 0 0 0 0 45 0 0 144 2
616 767
76 767
1 0 29 0 0 0 0 45 0 0 136 2
616 749
425 749
0 2 31 0 0 8320 0 0 41 75 0 5
1077 652
1077 1028
601 1028
601 936
616 936
3 0 9 0 0 0 0 37 0 0 0 2
1061 972
1184 972
4 2 32 0 0 12416 0 36 37 0 0 4
985 999
991 999
991 981
1015 981
3 1 33 0 0 4224 0 38 37 0 0 4
990 956
1008 956
1008 963
1015 963
0 3 34 0 0 8320 0 0 36 63 0 3
784 858
784 1008
940 1008
0 1 35 0 0 4224 0 0 36 64 0 3
826 793
826 990
940 990
0 2 36 0 0 8192 0 0 38 61 0 3
884 927
884 965
945 965
1 0 37 0 0 8320 0 38 0 0 62 3
945 947
926 947
926 825
3 2 36 0 0 4224 0 41 39 0 0 4
661 927
973 927
973 862
989 862
3 1 37 0 0 0 0 40 39 0 0 3
914 825
989 825
989 844
3 2 34 0 0 0 0 42 40 0 0 4
735 858
858 858
858 834
865 834
3 1 35 0 0 0 0 47 40 0 0 4
813 793
846 793
846 816
865 816
3 2 38 0 0 8320 0 43 42 0 0 3
660 883
660 867
689 867
3 1 39 0 0 8320 0 44 42 0 0 3
661 838
661 849
689 849
4 1 40 0 0 8320 0 46 47 0 0 3
736 782
736 784
767 784
3 1 41 0 0 4224 0 45 46 0 0 4
665 758
682 758
682 773
691 773
0 2 42 0 0 8320 0 0 54 95 0 5
1033 331
1033 708
557 708
557 616
572 616
2 0 43 0 0 4096 0 48 0 0 139 2
723 482
296 482
1 0 44 0 0 4096 0 52 0 0 123 2
571 554
500 554
1 0 45 0 0 4096 0 51 0 0 135 2
572 509
465 509
2 0 11 0 0 0 0 50 0 0 144 2
572 447
76 447
1 0 45 0 0 0 0 50 0 0 135 2
572 429
465 429
3 0 31 0 0 0 0 59 0 0 0 2
1017 652
1140 652
3 2 46 0 0 8320 0 58 59 0 0 3
947 679
947 661
971 661
3 1 47 0 0 4224 0 57 59 0 0 4
946 636
964 636
964 643
971 643
0 2 48 0 0 8320 0 0 58 84 0 3
740 538
740 688
902 688
0 1 49 0 0 4224 0 0 58 85 0 3
782 473
782 670
902 670
0 2 50 0 0 8192 0 0 57 82 0 3
840 607
840 645
901 645
1 0 51 0 0 8320 0 57 0 0 83 3
901 627
882 627
882 505
3 2 50 0 0 4224 0 54 56 0 0 4
617 607
929 607
929 542
945 542
3 1 51 0 0 0 0 55 56 0 0 3
870 505
945 505
945 524
3 2 48 0 0 0 0 53 55 0 0 4
691 538
814 538
814 514
821 514
3 1 49 0 0 0 0 48 55 0 0 4
769 473
802 473
802 496
821 496
1 0 10 0 0 0 0 54 0 0 127 2
572 598
70 598
3 2 52 0 0 8320 0 52 53 0 0 3
616 563
616 547
645 547
3 1 53 0 0 8320 0 51 53 0 0 3
617 518
617 529
645 529
2 0 11 0 0 0 0 52 0 0 144 2
571 572
76 572
2 0 13 0 0 0 0 51 0 0 143 2
572 527
121 527
4 1 54 0 0 8320 0 49 48 0 0 3
692 462
692 464
723 464
3 1 55 0 0 4224 0 50 49 0 0 4
621 438
638 438
638 453
647 453
2 0 17 0 0 0 0 49 0 0 126 2
647 462
156 462
3 0 16 0 0 0 0 49 0 0 145 2
647 471
35 471
3 0 42 0 0 0 0 60 0 0 0 2
1018 331
1141 331
3 1 6 0 0 4224 0 63 19 0 0 3
995 212
1362 212
1362 60
3 2 56 0 0 8320 0 61 60 0 0 3
948 358
948 340
972 340
3 1 57 0 0 4224 0 62 60 0 0 4
947 315
965 315
965 322
972 322
0 2 58 0 0 8320 0 0 61 105 0 3
741 217
741 367
903 367
0 1 59 0 0 4224 0 0 61 106 0 3
783 152
783 349
903 349
0 2 60 0 0 8192 0 0 62 103 0 3
841 286
841 324
902 324
1 0 61 0 0 8320 0 62 0 0 104 3
902 306
883 306
883 184
3 2 60 0 0 4224 0 65 63 0 0 4
618 286
930 286
930 221
946 221
3 1 61 0 0 0 0 64 63 0 0 3
871 184
946 184
946 203
3 2 58 0 0 0 0 66 64 0 0 4
692 217
815 217
815 193
822 193
3 1 59 0 0 0 0 77 64 0 0 4
770 152
803 152
803 175
822 175
2 0 62 0 0 4096 0 65 0 0 142 2
573 295
170 295
1 0 10 0 0 0 0 65 0 0 127 2
573 277
70 277
3 2 63 0 0 8320 0 67 66 0 0 3
617 242
617 226
646 226
3 1 64 0 0 8320 0 68 66 0 0 3
618 197
618 208
646 208
2 0 11 0 0 0 0 67 0 0 144 2
572 251
76 251
1 0 65 0 0 4096 0 67 0 0 122 2
572 233
542 233
2 0 13 0 0 0 0 68 0 0 143 2
573 206
121 206
1 0 66 0 0 4096 0 68 0 0 134 2
573 188
508 188
2 0 67 0 0 4096 0 77 0 0 138 2
724 161
336 161
4 1 68 0 0 8320 0 76 77 0 0 3
693 141
693 143
724 143
3 1 69 0 0 4224 0 75 76 0 0 4
622 117
639 117
639 132
648 132
2 0 17 0 0 0 0 76 0 0 126 2
648 141
156 141
3 0 16 0 0 0 0 76 0 0 145 2
648 150
35 150
2 0 11 0 0 0 0 75 0 0 144 2
573 126
76 126
1 0 66 0 0 0 0 75 0 0 134 2
573 108
508 108
2 0 65 0 0 4224 0 69 0 0 0 2
542 78
542 1533
2 0 44 0 0 4224 0 70 0 0 0 2
500 77
500 1528
2 0 28 0 0 4224 0 71 0 0 0 2
460 77
460 1527
2 0 12 0 0 4224 0 72 0 0 0 2
418 78
418 1524
2 0 17 0 0 4224 0 73 0 0 0 2
156 73
156 1526
2 0 10 0 0 4224 0 74 0 0 0 2
70 74
70 1526
1 0 66 0 0 0 0 69 0 0 134 2
506 78
508 78
1 0 45 0 0 0 0 70 0 0 135 2
464 77
465 77
1 0 29 0 0 0 0 71 0 0 136 2
424 77
425 77
1 0 14 0 0 0 0 72 0 0 137 2
382 78
381 78
1 0 13 0 0 0 0 73 0 0 143 2
120 73
121 73
1 0 16 0 0 0 0 74 0 0 145 2
34 74
35 74
1 0 66 0 0 4224 0 1 0 0 0 2
508 65
508 1531
1 0 45 0 0 4224 0 2 0 0 0 2
465 64
465 1525
1 0 29 0 0 4224 0 3 0 0 0 2
425 64
425 1524
1 0 14 0 0 4224 0 4 0 0 0 2
381 66
381 1522
1 0 67 0 0 4224 0 5 0 0 0 2
336 65
336 1525
1 0 43 0 0 4224 0 6 0 0 0 2
296 66
296 1525
1 0 30 0 0 4224 0 7 0 0 0 2
252 68
252 1525
1 0 15 0 0 4224 0 8 0 0 0 2
214 65
214 1527
1 0 62 0 0 4224 0 9 0 0 0 2
170 67
170 1526
1 0 13 0 0 4224 0 10 0 0 0 2
121 67
121 1527
1 0 11 0 0 4224 0 11 0 0 0 2
76 67
76 1527
1 0 16 0 0 4224 0 12 0 0 0 2
35 68
35 1526
54
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 8
604 29 693 60
611 33 685 54
8 56 gates
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1698 4 1727 35
1705 8 1719 29
1 C
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1635 3 1662 34
1642 7 1654 28
1 S
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1542 8 1571 39
1549 12 1563 33
1 Z
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1431 7 1459 38
1438 11 1451 32
1 V
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1132 -1 1173 30
1139 3 1165 24
2 C5
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1190 -2 1231 29
1197 2 1223 23
2 F4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1242 -2 1283 29
1249 2 1275 23
2 F3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1300 -1 1342 30
1307 3 1334 24
2 F2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1065 1256 1106 1287
1072 1260 1098 1281
2 C5
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1035 1126 1076 1157
1042 1130 1068 1151
2 F4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
686 1215 727 1246
693 1219 719 1240
2 Z4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
735 1136 775 1167
742 1140 767 1161
2 Y4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
791 1058 831 1089
798 1062 823 1083
2 X4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1052 936 1093 967
1059 940 1085 961
2 C4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1022 806 1063 837
1029 810 1055 831
2 F3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
673 895 714 926
680 899 706 920
2 Z3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
722 816 762 847
729 820 754 841
2 Y3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
778 738 818 769
785 742 810 763
2 X3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
978 486 1020 517
985 490 1012 511
2 F2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1008 616 1049 647
1015 620 1041 641
2 C3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
629 575 671 606
636 579 663 600
2 Z2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
678 496 719 527
685 500 711 521
2 Y2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
734 418 775 449
741 422 767 443
2 X2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1004 276 1046 307
1011 280 1038 301
2 C2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
1349 0 1381 31
1353 4 1376 25
2 F1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
983 159 1015 190
987 163 1010 184
2 F1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
620 250 652 281
624 254 647 275
2 Z1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
692 176 723 207
696 180 718 201
2 Y1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
763 105 794 136
767 109 789 130
2 X1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
32 975 67 1006
38 979 60 1000
2 s2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
62 977 89 1008
66 981 84 1002
2 s1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
124 969 155 1000
128 973 150 994
2 s0
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
160 979 192 1010
164 983 187 1004
2 C1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
198 977 232 1008
202 981 227 1002
2 A4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
234 981 268 1012
238 985 263 1006
2 A3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
278 980 313 1011
282 984 308 1005
2 A2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
322 978 353 1009
326 982 348 1003
2 A1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
383 959 419 990
387 963 414 984
2 B4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
426 962 462 993
430 966 457 987
2 B3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
509 962 542 993
513 966 537 987
2 B1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
462 952 505 1009
469 956 497 998
2 B2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
449 -2 492 55
456 2 484 44
2 B2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
492 -1 525 30
496 3 520 24
2 B1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
408 -2 444 29
412 2 439 23
2 B3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
367 -2 403 29
371 2 398 23
2 B4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
321 -4 352 27
325 0 347 21
2 A1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
280 -4 315 27
284 0 310 21
2 A2
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
238 -3 272 28
242 1 267 22
2 A3
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
199 -4 233 27
203 0 228 21
2 A4
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
156 -4 188 27
160 0 183 21
2 C1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
105 -4 136 27
109 0 131 21
2 s0
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
62 -4 89 27
66 0 84 21
2 s1
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 2
21 -2 56 29
27 2 49 23
2 s2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
