CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
3
7 Ground~
168 241 69 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
42655.5 0
0
7 74LS173
129 141 78 0 1 29
0 0
0
0 0 4832 0
7 74LS173
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
391 0 0
2
42655.4 0
0
7 74LS173
129 335 62 0 1 29
0 0
0
0 0 4832 0
7 74LS173
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
3124 0 0
2
42655.4 0
0
33
1 0 0 0 0 0 0 3 0 0 6 3
303 35
241 35
241 56
0 0 0 0 0 0 0 0 0 3 0 5
257 360
753 360
753 193
772 193
772 209
4 4 0 0 0 0 0 3 2 0 0 6
303 62
257 62
257 361
13 361
13 78
109 78
0 0 0 0 0 0 0 0 0 5 0 5
373 39
389 39
389 12
705 12
705 145
10 9 0 0 0 0 0 3 3 0 0 2
373 44
373 35
0 1 0 0 0 0 0 0 1 7 0 3
179 56
241 56
241 63
10 9 0 0 0 0 0 2 2 0 0 2
179 60
179 51
0 0 0 0 0 0 0 0 0 10 9 6
297 49
290 49
290 6
597 6
597 111
659 111
0 0 0 0 0 0 0 0 0 11 0 5
103 63
39 63
39 341
659 341
659 83
3 2 0 0 0 0 0 3 3 0 0 2
297 53
297 44
3 2 0 0 0 0 0 2 2 0 0 2
103 69
103 60
6 0 0 0 0 0 0 2 0 0 25 5
109 96
77 96
77 282
429 282
429 275
7 0 0 0 0 0 0 2 0 0 30 4
109 105
94 105
94 268
447 268
8 0 0 0 0 0 0 2 0 0 26 3
109 114
109 256
470 256
5 0 0 0 0 0 0 3 0 0 33 4
303 71
267 71
267 245
491 245
6 0 0 0 0 0 0 3 0 0 27 4
303 80
297 80
297 228
514 228
7 0 0 0 0 0 0 3 0 0 31 4
303 89
278 89
278 206
537 206
8 0 0 0 0 0 0 3 0 0 28 4
303 98
303 193
560 193
560 118
11 0 0 0 0 0 0 2 0 0 29 4
173 87
287 87
287 137
411 137
12 0 0 0 0 0 0 2 0 0 25 4
173 96
283 96
283 146
429 146
13 0 0 0 0 0 0 2 0 0 30 4
173 105
272 105
272 156
447 156
14 0 0 0 0 0 0 2 0 0 26 4
173 114
218 114
218 173
470 173
12 0 0 0 0 0 0 3 0 0 27 4
367 80
499 80
499 100
514 100
13 0 0 0 0 0 0 3 0 0 31 4
367 89
522 89
522 109
537 109
0 0 0 0 0 0 0 0 0 0 0 2
429 279
429 49
0 0 0 0 0 0 0 0 0 0 0 2
470 280
470 49
0 0 0 0 0 0 0 0 0 0 0 2
514 280
514 49
14 0 0 0 0 0 0 3 0 0 0 5
367 98
560 98
560 118
560 118
560 49
0 5 0 0 0 0 0 0 2 0 0 5
411 49
411 310
56 310
56 87
109 87
0 0 0 0 0 0 0 0 0 0 0 2
447 48
447 280
0 0 0 0 0 0 0 0 0 0 0 2
537 49
537 281
11 0 0 0 0 0 0 3 0 0 0 3
367 71
491 71
491 49
0 0 0 0 0 0 0 0 0 32 0 2
491 53
491 280
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
77 37 116 61
84 42 108 58
3 CLR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
769 217 808 241
776 223 800 239
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
703 153 742 177
710 158 734 174
3 Ei'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
643 41 682 65
650 46 674 62
3 Li'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
395 25 422 49
400 29 416 45
2 I7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
415 23 442 47
420 27 436 43
2 I6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
437 24 464 48
442 28 458 44
2 I5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
462 25 489 49
467 29 483 45
2 I4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
482 25 509 49
487 29 503 45
2 I3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
503 25 530 49
508 29 524 45
2 I2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
525 25 552 49
530 29 546 45
2 I1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
548 24 575 48
553 28 569 44
2 I0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
100 7 271 31
105 11 265 27
20 INSTRUCTION REGISTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
467 10 518 34
472 14 512 30
5 W BUS
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
