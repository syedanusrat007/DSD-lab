CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
940 420 15 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
111
13 Logic Switch~
5 445 1602 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5267 0 0
2
42987.8 0
0
13 Logic Switch~
5 206 441 0 10 11
0 74 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8838 0 0
2
42987.8 0
0
13 Logic Switch~
5 380 501 0 10 11
0 75 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V20
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7159 0 0
2
5.89815e-315 5.30499e-315
0
13 Logic Switch~
5 348 500 0 1 11
0 76
0
0 0 21360 90
2 0V
11 0 25 8
3 V22
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5812 0 0
2
5.89815e-315 5.32571e-315
0
13 Logic Switch~
5 317 500 0 10 11
0 77 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V23
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
331 0 0
2
5.89815e-315 5.34643e-315
0
13 Logic Switch~
5 284 498 0 10 11
0 78 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V24
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9604 0 0
2
5.89815e-315 5.3568e-315
0
13 Logic Switch~
5 1536 965 0 1 11
0 97
0
0 0 21360 90
2 0V
11 0 25 8
3 V12
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7518 0 0
2
5.89815e-315 5.36716e-315
0
13 Logic Switch~
5 1569 967 0 1 11
0 96
0
0 0 21360 90
2 0V
11 0 25 8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4832 0 0
2
5.89815e-315 5.37752e-315
0
13 Logic Switch~
5 1600 967 0 1 11
0 95
0
0 0 21360 90
2 0V
11 0 25 8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6798 0 0
2
5.89815e-315 5.38788e-315
0
13 Logic Switch~
5 1632 968 0 10 11
0 94 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3336 0 0
2
5.89815e-315 5.39306e-315
0
13 Logic Switch~
5 1385 966 0 10 11
0 86 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8370 0 0
2
5.89815e-315 5.39824e-315
0
13 Logic Switch~
5 1353 965 0 1 11
0 85
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3910 0 0
2
5.89815e-315 5.40342e-315
0
13 Logic Switch~
5 1322 965 0 1 11
0 84
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
316 0 0
2
5.89815e-315 5.4086e-315
0
13 Logic Switch~
5 1289 963 0 1 11
0 83
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
536 0 0
2
5.89815e-315 5.41378e-315
0
7 74LS125
115 850 1176 0 12 25
0 4 87 4 88 4 89 4 3 8
7 6 5
0
0 0 4848 0
7 74LS125
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 0 0 0 0
1 U
4460 0 0
2
42987.9 0
0
7 74LS125
115 1102 852 0 12 25
0 9 83 9 84 9 85 9 86 5
6 7 8
0
0 0 4848 180
7 74LS125
-24 -51 25 -43
2 U4
-13 -52 1 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 0 0 0 0
1 U
3260 0 0
2
42987.9 0
0
7 74LS125
115 1091 430 0 12 25
0 10 62 10 63 10 64 10 65 5
6 7 8
0
0 0 4848 180
7 74LS125
-24 -51 25 -43
3 U15
-16 -52 5 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 0 0 0 0
1 U
5156 0 0
2
42987.9 0
0
7 74LS125
115 1098 294 0 12 25
0 11 58 11 59 11 60 11 61 5
6 7 8
0
0 0 4848 180
7 74LS125
-24 -51 25 -43
2 U2
-13 -52 1 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 0 0 0 0
1 U
3133 0 0
2
42987.9 0
0
7 74LS125
115 829 169 0 12 25
0 12 82 12 81 12 13 12 80 5
6 7 8
0
0 0 4848 0
7 74LS125
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 0 0 0 0
1 U
5523 0 0
2
42987.9 0
0
14 Logic Display~
6 1708 2107 0 1 2
10 16
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L48
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3746 0 0
2
5.89815e-315 0
0
5 4049~
219 1698 1918 0 2 22
0 11 16
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U26D
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 9 0
1 U
5668 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1625 2100 0 1 2
10 9
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L47
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5368 0 0
2
5.89815e-315 0
0
5 4049~
219 1861 705 0 2 22
0 18 17
0
0 0 624 180
4 4049
-7 -24 21 -16
4 U26C
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 9 0
1 U
8293 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1505 2028 0 1 2
10 21
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L46
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3232 0 0
2
5.89815e-315 0
0
5 4071~
219 1504 1658 0 3 22
0 18 20 21
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U30B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 13 0
1 U
6644 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1439 2027 0 1 2
10 15
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L45
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4978 0 0
2
5.89815e-315 0
0
5 4071~
219 1436 1658 0 3 22
0 19 18 15
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U30A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
9207 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1365 2019 0 1 2
10 10
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L44
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6998 0 0
2
5.89815e-315 0
0
9 2-In AND~
219 1368 1706 0 3 22
0 15 9 10
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U28B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3175 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1316 2002 0 1 2
10 11
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L43
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3378 0 0
2
5.89815e-315 0
0
9 2-In AND~
219 1318 1740 0 3 22
0 9 22 11
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U28A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
922 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1230 1981 0 1 2
10 23
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L42
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6891 0 0
2
5.89815e-315 0
0
5 4001~
219 1225 1775 0 3 22
0 25 24 23
0
0 0 624 270
4 4001
-14 -24 14 -16
4 U25C
32 -10 60 -2
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 8 0
1 U
5407 0 0
2
5.89815e-315 0
0
9 2-In AND~
219 1241 1713 0 3 22
0 26 9 25
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7349 0 0
2
5.89815e-315 0
0
8 4-In OR~
219 1246 1646 0 5 22
0 19 18 98 27 26
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U27A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 10 0
1 U
3919 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1162 1973 0 1 2
10 4
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L41
19 -2 40 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9747 0 0
2
5.89815e-315 0
0
5 4049~
219 1161 1808 0 2 22
0 28 4
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U26B
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 9 0
1 U
5310 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 1119 1978 0 1 2
10 29
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4318 0 0
2
5.89815e-315 0
0
5 4049~
219 1116 1810 0 2 22
0 30 29
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U26A
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 9 0
1 U
3917 0 0
2
5.89815e-315 0
0
5 4001~
219 1055 1715 0 3 22
0 24 30 31
0
0 0 624 270
4 4001
-14 -24 14 -16
4 U25B
32 -10 60 -2
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 8 0
1 U
7930 0 0
2
5.89815e-315 0
0
5 4001~
219 960 1713 0 3 22
0 28 12 32
0
0 0 624 270
4 4001
-14 -24 14 -16
4 U25A
32 -10 60 -2
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 8 0
1 U
6128 0 0
2
5.89815e-315 0
0
9 2-In AND~
219 1072 1659 0 3 22
0 34 33 24
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7346 0 0
2
5.89815e-315 5.32571e-315
0
14 Logic Display~
6 1052 1982 0 1 2
10 31
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L39
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8577 0 0
2
5.89815e-315 0
0
9 2-In AND~
219 977 1655 0 3 22
0 33 9 28
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3372 0 0
2
5.89815e-315 5.32571e-315
0
14 Logic Display~
6 955 1978 0 1 2
10 32
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L38
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3741 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 876 1962 0 1 2
10 35
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L37
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5813 0 0
2
5.89815e-315 0
0
5 4011~
219 877 1784 0 3 22
0 36 9 35
0
0 0 624 270
4 4011
-7 -24 21 -16
4 U24A
20 -7 48 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 7 0
1 U
3213 0 0
2
5.89815e-315 0
0
8 2-In OR~
219 885 1716 0 3 22
0 38 37 36
0
0 0 624 270
5 74F32
-18 -24 17 -16
4 U23A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3694 0 0
2
5.89815e-315 0
0
9 2-In AND~
219 899 1660 0 3 22
0 39 40 38
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U22A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4327 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 826 1956 0 1 2
10 30
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L36
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8800 0 0
2
5.89815e-315 0
0
14 Logic Display~
6 793 1962 0 1 2
10 12
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L35
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3406 0 0
2
5.89815e-315 0
0
9 2-In XOR~
219 386 1369 0 3 22
0 2 12 41
0
0 0 624 90
6 74LS86
-21 -24 21 -16
4 U31A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
6455 0 0
2
5.89815e-315 5.41896e-315
0
7 Ground~
168 380 1392 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9319 0 0
2
5.89815e-315 5.42414e-315
0
7 Ground~
168 571 1263 0 1 3
0 2
0
0 0 53360 180
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3172 0 0
2
5.89815e-315 5.42933e-315
0
2 +V
167 675 1372 0 1 3
0 54
0
0 0 54256 180
3 10V
6 -2 27 6
3 V32
6 -12 27 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
38 0 0
2
42987.8 3
0
9 3-In NOR~
219 711 1261 0 4 22
0 12 30 9 55
0
0 0 624 180
5 74F27
-18 -24 17 -16
4 U21A
-11 -2 17 6
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
376 0 0
2
42987.8 4
0
14 Logic Display~
6 1552 1300 0 1 2
10 9
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L33
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6666 0 0
2
42987.8 5
0
14 Logic Display~
6 1552 1325 0 1 2
10 30
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L32
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9365 0 0
2
42987.8 6
0
14 Logic Display~
6 1552 1351 0 1 2
10 12
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L31
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3251 0 0
2
42987.8 7
0
14 Logic Display~
6 1552 1274 0 1 2
10 34
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L30
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5481 0 0
2
42987.8 8
0
7 74LS164
127 716 1324 0 12 25
0 55 55 14 54 99 100 101 102 34
9 30 12
0
0 0 4848 0
6 74F164
-21 -51 21 -43
3 U20
-14 4 7 12
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
7788 0 0
2
42987.8 9
0
14 Logic Display~
6 1702 1406 0 1 2
10 33
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L21
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3273 0 0
2
5.89815e-315 5.44487e-315
0
14 Logic Display~
6 1700 1481 0 1 2
10 20
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L23
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3761 0 0
2
5.89815e-315 5.44746e-315
0
14 Logic Display~
6 1700 1455 0 1 2
10 18
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L24
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
5.89815e-315 5.45005e-315
0
14 Logic Display~
6 1695 1556 0 1 2
10 37
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L25
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4244 0 0
2
5.89815e-315 5.45264e-315
0
14 Logic Display~
6 1693 1579 0 1 2
10 40
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L26
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5225 0 0
2
5.89815e-315 5.45523e-315
0
14 Logic Display~
6 1697 1534 0 1 2
10 22
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L27
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
768 0 0
2
5.89815e-315 5.45782e-315
0
14 Logic Display~
6 1698 1505 0 1 2
10 27
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L28
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5735 0 0
2
5.89815e-315 5.46041e-315
0
14 Logic Display~
6 1693 1608 0 1 2
10 56
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L29
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5881 0 0
2
5.89815e-315 5.463e-315
0
14 Logic Display~
6 1701 1431 0 1 2
10 19
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3275 0 0
2
5.89815e-315 5.46559e-315
0
7 74LS154
95 551 1316 0 22 45
0 2 2 50 51 52 53 103 104 105
106 107 108 56 40 37 22 27 20 18
19 33 109
0
0 0 4848 270
6 74F154
-21 -87 21 -79
3 U17
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
4203 0 0
2
5.89815e-315 5.48113e-315
0
9 4-In NOR~
219 1422 275 0 5 22
0 61 60 59 58 39
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 1 0
1 U
3440 0 0
2
5.89815e-315 5.48243e-315
0
7 74LS181
132 1190 471 0 22 45
0 15 20 21 15 58 59 60 61 69
68 67 66 19 18 110 111 112 113 62
63 64 65
0
0 0 4848 180
7 74LS181
-24 -69 25 -61
3 U14
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
9102 0 0
2
5.89815e-315 5.48631e-315
0
6 PROM32
80 777 600 0 14 29
0 31 2 45 44 43 42 49 48 47
46 5 6 7 8
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5586 0 0
2
5.89815e-315 5.48761e-315
0
DAJAAAAAAAAAAAAAAAAAAFAAAAAAAAAFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 Ground~
168 389 599 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
525 0 0
2
5.89815e-315 5.4889e-315
0
7 74LS173
129 771 440 0 14 29
0 2 32 32 14 8 7 6 5 2
2 70 71 72 73
0
0 0 4848 270
6 74F173
-21 -51 21 -43
3 U12
47 -2 68 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6206 0 0
2
5.89815e-315 5.4902e-315
0
7 Ground~
168 869 405 0 1 3
0 2
0
0 0 53360 90
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3418 0 0
2
5.89815e-315 5.49149e-315
0
7 Ground~
168 546 479 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9312 0 0
2
5.89815e-315 5.49279e-315
0
7 74LS257
147 614 517 0 14 29
0 74 70 75 71 76 72 77 73 78
2 42 43 44 45
0
0 0 4848 270
6 74F257
-21 -60 21 -52
3 U11
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
7419 0 0
2
5.89815e-315 5.49408e-315
0
7 Ground~
168 475 168 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
472 0 0
2
5.89815e-315 5.49538e-315
0
2 +V
167 598 114 0 1 3
0 79
0
0 0 54256 0
2 5V
-8 -22 6 -14
3 V17
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4714 0 0
2
5.89815e-315 5.49667e-315
0
7 74LS193
137 663 168 0 14 29
0 30 79 35 2 5 6 7 8 114
115 82 81 13 80
0
0 0 4848 0
6 74F193
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9386 0 0
2
5.89815e-315 5.49797e-315
0
7 Ground~
168 743 1174 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7610 0 0
2
5.89815e-315 5.50185e-315
0
7 74LS173
129 671 1128 0 14 29
0 2 29 29 14 8 7 6 5 2
2 87 88 89 3
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U7
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3482 0 0
2
5.89815e-315 5.50315e-315
0
7 74LS173
129 542 1127 0 14 29
0 41 29 29 14 46 47 48 49 2
2 53 52 51 50
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U6
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3608 0 0
2
5.89815e-315 5.50444e-315
0
14 Logic Display~
6 1390 1160 0 1 2
10 93
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6397 0 0
2
5.89815e-315 5.50574e-315
0
14 Logic Display~
6 1370 1160 0 1 2
10 92
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3967 0 0
2
5.89815e-315 5.50703e-315
0
14 Logic Display~
6 1350 1160 0 1 2
10 91
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8621 0 0
2
5.89815e-315 5.50833e-315
0
14 Logic Display~
6 1331 1160 0 1 2
10 90
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89815e-315 5.50963e-315
0
7 Ground~
168 1253 1131 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7385 0 0
2
5.89815e-315 5.51092e-315
0
7 74LS173
129 1158 1090 0 14 29
0 2 16 16 14 5 6 7 8 2
2 90 91 92 93
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U5
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6519 0 0
2
5.89815e-315 5.51222e-315
0
7 Ground~
168 1400 746 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
552 0 0
2
5.89815e-315 5.51286e-315
0
7 74LS257
147 1323 708 0 14 29
0 17 83 97 84 96 85 95 86 94
2 69 68 67 66
0
0 0 4848 90
6 74F257
-21 -60 21 -52
2 U3
54 -6 68 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
5551 0 0
2
5.89815e-315 5.51416e-315
0
7 Ground~
168 1254 242 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8715 0 0
2
5.89815e-315 5.51545e-315
0
7 74LS173
129 1159 200 0 14 29
0 2 23 23 14 5 6 7 8 2
2 58 59 60 61
0
0 0 4848 270
6 74F173
-21 -51 21 -43
2 U1
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
9763 0 0
2
5.89815e-315 5.5161e-315
0
14 Logic Display~
6 916 1239 0 1 2
10 49
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L16
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8443 0 0
2
42987.8 10
0
14 Logic Display~
6 935 1239 0 1 2
10 48
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L15
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3719 0 0
2
42987.8 11
0
14 Logic Display~
6 955 1239 0 1 2
10 47
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L14
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8671 0 0
2
42987.8 12
0
14 Logic Display~
6 975 1239 0 1 2
10 46
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L13
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
42987.8 13
0
14 Logic Display~
6 1053 1239 0 1 2
10 8
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L12
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
49 0 0
2
42987.8 14
0
14 Logic Display~
6 1033 1239 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L11
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6536 0 0
2
42987.8 15
0
14 Logic Display~
6 1013 1239 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L10
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3931 0 0
2
42987.8 16
0
14 Logic Display~
6 994 1239 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4390 0 0
2
42987.8 17
0
14 Logic Display~
6 994 94 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3242 0 0
2
42987.8 18
0
14 Logic Display~
6 1013 94 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6760 0 0
2
42987.8 19
0
14 Logic Display~
6 1033 94 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5760 0 0
2
42987.8 20
0
14 Logic Display~
6 1053 94 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3781 0 0
2
42987.8 21
0
14 Logic Display~
6 975 94 0 1 2
10 46
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8545 0 0
2
42987.8 22
0
14 Logic Display~
6 955 94 0 1 2
10 47
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9739 0 0
2
42987.8 23
0
14 Logic Display~
6 935 94 0 1 2
10 48
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
388 0 0
2
42987.8 24
0
14 Logic Display~
6 916 94 0 1 2
10 49
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
42987.8 25
0
286
0 8 3 0 0 4096 0 0 15 232 0 2
810 1212
818 1212
5 0 4 0 0 12288 0 15 0 0 4 4
812 1185
799 1185
799 1178
775 1178
3 0 4 0 0 4096 0 15 0 0 4 2
812 1167
775 1167
1 0 4 0 0 8192 0 15 0 0 224 3
812 1149
775 1149
775 1203
12 0 5 0 0 0 0 15 0 0 226 2
882 1212
882 1212
11 0 6 0 0 0 0 15 0 0 227 2
882 1194
882 1194
10 0 7 0 0 0 0 15 0 0 228 2
882 1176
882 1176
9 0 8 0 0 0 0 15 0 0 229 2
882 1158
882 1158
7 0 9 0 0 0 0 16 0 0 43 2
1134 829
1134 829
5 0 9 0 0 0 0 16 0 0 42 2
1134 847
1134 847
3 0 9 0 0 0 0 16 0 0 41 2
1134 865
1134 865
1 0 9 0 0 0 0 16 0 0 46 2
1134 883
1134 883
12 0 8 0 0 0 0 17 0 0 279 2
1053 398
1053 398
11 0 7 0 0 0 0 17 0 0 180 2
1053 416
1053 416
10 0 6 0 0 0 0 17 0 0 179 2
1053 434
1053 434
9 0 5 0 0 0 0 17 0 0 178 2
1053 452
1053 452
7 0 10 0 0 4096 0 17 0 0 63 2
1123 407
1126 407
5 0 10 0 0 0 0 17 0 0 63 2
1123 425
1126 425
3 0 10 0 0 0 0 17 0 0 63 2
1123 443
1126 443
1 0 10 0 0 0 0 17 0 0 63 2
1123 461
1126 461
1 0 11 0 0 4096 0 18 0 0 24 2
1130 325
1168 325
3 0 11 0 0 0 0 18 0 0 24 2
1130 307
1168 307
5 0 11 0 0 0 0 18 0 0 24 2
1130 289
1168 289
7 0 11 0 0 8192 0 18 0 0 25 3
1130 271
1168 271
1168 340
0 0 11 0 0 8320 0 0 0 68 0 4
1316 1848
2081 1848
2081 340
1144 340
5 0 12 0 0 4096 0 19 0 0 29 2
791 178
775 178
3 0 12 0 0 0 0 19 0 0 29 2
791 160
775 160
1 0 12 0 0 0 0 19 0 0 29 2
791 142
775 142
7 0 12 0 0 16512 0 19 0 0 116 6
791 196
775 196
775 100
57 100
57 1809
793 1809
6 0 13 0 0 4096 0 19 0 0 217 2
797 187
789 187
12 0 8 0 0 0 0 19 0 0 209 2
861 205
861 205
11 0 7 0 0 0 0 19 0 0 208 2
861 187
861 187
10 0 6 0 0 0 0 19 0 0 207 2
861 169
861 169
9 0 5 0 0 0 0 19 0 0 206 2
861 151
861 151
1 0 14 0 0 12304 0 1 0 0 117 4
457 1602
457 1484
345 1484
345 1234
1 0 15 0 0 12288 0 29 0 0 60 5
1375 1684
1375 1666
1410 1666
1410 1718
1446 1718
2 0 16 0 0 4096 0 91 0 0 38 2
1178 1054
1178 1012
3 0 16 0 0 12416 0 91 0 0 39 5
1169 1054
1169 1012
1962 1012
1962 1966
1705 1966
1 2 16 0 0 0 0 20 21 0 0 6
1708 2093
1705 2093
1705 1943
1700 1943
1700 1936
1701 1936
0 1 11 0 0 0 0 0 21 68 0 3
1316 1799
1701 1799
1701 1900
0 0 9 0 0 4096 0 0 0 0 44 2
1127 865
1141 865
0 0 9 0 0 0 0 0 0 0 44 2
1127 847
1141 847
0 0 9 0 0 0 0 0 0 0 44 2
1127 829
1141 829
0 0 9 0 0 8320 0 0 0 45 46 5
1632 1781
1978 1781
1978 803
1141 803
1141 883
1 0 9 0 0 0 0 22 0 0 149 9
1625 2086
1632 2086
1632 1761
1628 1761
1628 1728
1637 1728
1637 1376
1416 1376
1416 1304
0 0 9 0 0 0 0 0 0 0 0 2
1127 883
1146 883
4 0 14 0 0 8192 0 91 0 0 118 3
1160 1060
1160 1037
2152 1037
2 1 17 0 0 4224 0 23 93 0 0 5
1846 705
1453 705
1453 767
1282 767
1282 739
1 0 18 0 0 4096 0 23 0 0 51 2
1882 705
2011 705
0 13 19 0 0 12416 0 0 73 159 0 7
1587 1435
1587 1710
1997 1710
1997 560
1142 560
1142 520
1158 520
14 0 18 0 0 16512 0 73 0 0 158 7
1158 511
1134 511
1134 542
2011 542
2011 1676
1570 1676
1570 1459
2 0 20 0 0 8320 0 73 0 0 157 5
1222 511
2026 511
2026 1650
1548 1650
1548 1485
0 3 21 0 0 8320 0 0 73 54 0 4
1512 1862
2053 1862
2053 502
1222 502
1 3 21 0 0 0 0 24 25 0 0 5
1505 2014
1512 2014
1512 1689
1507 1689
1507 1688
2 0 20 0 0 0 0 25 0 0 157 2
1498 1642
1498 1485
1 0 18 0 0 0 0 25 0 0 158 2
1516 1642
1516 1459
1 0 15 0 0 4096 0 73 0 0 59 3
1222 520
1410 520
1410 493
0 0 15 0 0 4096 0 0 0 59 60 2
2037 1872
1446 1872
4 0 15 0 0 8320 0 73 0 0 0 3
1222 493
2037 493
2037 1876
1 3 15 0 0 0 0 26 27 0 0 4
1439 2013
1446 2013
1446 1688
1439 1688
2 0 18 0 0 0 0 27 0 0 158 4
1430 1642
1430 1475
1431 1475
1431 1460
1 0 19 0 0 0 0 27 0 0 159 4
1448 1642
1448 1450
1449 1450
1449 1435
0 0 10 0 0 8320 0 0 0 65 0 6
1365 1839
2067 1839
2067 369
1126 369
1126 461
1121 461
2 0 9 0 0 0 0 29 0 0 149 2
1357 1684
1357 1304
1 3 10 0 0 0 0 28 29 0 0 4
1365 2005
1365 1744
1366 1744
1366 1729
2 0 22 0 0 4096 0 31 0 0 155 2
1307 1718
1307 1537
1 0 9 0 0 0 0 31 0 0 149 2
1325 1718
1325 1304
1 3 11 0 0 0 0 30 31 0 0 2
1316 1988
1316 1763
2 0 23 0 0 4096 0 95 0 0 70 3
1179 164
1179 151
1170 151
3 0 23 0 0 12416 0 95 0 0 71 5
1170 164
1170 130
2102 130
2102 1819
1231 1819
1 3 23 0 0 0 0 32 33 0 0 3
1230 1967
1231 1967
1231 1808
0 2 24 0 0 4224 0 0 33 102 0 3
1070 1692
1222 1692
1222 1756
1 3 25 0 0 8320 0 33 34 0 0 3
1240 1756
1239 1756
1239 1736
2 0 9 0 0 0 0 34 0 0 149 2
1230 1691
1230 1304
5 1 26 0 0 8320 0 35 34 0 0 3
1249 1676
1248 1676
1248 1691
4 0 27 0 0 4096 0 35 0 0 156 2
1235 1626
1235 1511
2 0 18 0 0 0 0 35 0 0 158 2
1253 1626
1253 1460
1 0 19 0 0 0 0 35 0 0 159 2
1262 1626
1262 1435
4 0 14 0 0 0 0 95 0 0 118 3
1161 170
1161 109
2152 109
1 2 4 0 0 8192 0 36 37 0 0 4
1162 1959
1163 1959
1163 1826
1164 1826
0 1 28 0 0 4224 0 0 37 104 0 3
975 1683
1164 1683
1164 1790
3 0 29 0 0 4096 0 84 0 0 85 2
682 1092
682 1011
3 0 29 0 0 0 0 85 0 0 85 2
553 1091
553 1011
2 0 29 0 0 0 0 85 0 0 85 2
562 1091
562 1011
0 2 29 0 0 4224 0 0 84 86 0 5
1120 1851
13 1851
13 1011
691 1011
691 1092
2 1 29 0 0 0 0 39 38 0 0 4
1119 1828
1120 1828
1120 1964
1119 1964
0 1 30 0 0 4096 0 0 39 115 0 3
826 1630
1119 1630
1119 1792
4 0 14 0 0 0 0 84 0 0 89 3
673 1098
673 1031
544 1031
4 0 14 0 0 0 0 85 0 0 117 3
544 1097
544 1023
44 1023
1 0 31 0 0 8320 0 74 0 0 101 4
739 564
29 564
29 1836
1051 1836
4 0 14 0 0 0 0 76 0 0 117 3
773 410
773 299
44 299
3 0 32 0 0 4096 0 76 0 0 93 3
782 404
782 381
791 381
0 2 32 0 0 8320 0 0 76 103 0 5
956 1821
40 1821
40 287
791 287
791 404
2 0 30 0 0 4096 0 40 0 0 150 2
1052 1696
1052 1329
2 0 33 0 0 4096 0 42 0 0 160 2
1061 1637
1061 1409
1 0 34 0 0 4096 0 42 0 0 148 2
1079 1637
1079 1278
0 3 31 0 0 0 0 0 40 101 0 4
1051 1813
1051 1766
1061 1766
1061 1748
2 0 12 0 0 0 0 41 0 0 151 2
957 1694
957 1355
1 0 33 0 0 0 0 44 0 0 160 2
984 1633
984 1409
2 0 9 0 0 0 0 44 0 0 149 2
966 1633
966 1304
0 1 31 0 0 0 0 0 43 0 0 3
1051 1809
1051 1968
1052 1968
3 1 24 0 0 0 0 42 40 0 0 2
1070 1682
1070 1696
3 1 32 0 0 0 0 41 45 0 0 5
966 1746
966 1790
956 1790
956 1964
955 1964
3 1 28 0 0 0 0 44 41 0 0 2
975 1678
975 1694
0 3 35 0 0 8320 0 0 82 106 0 4
878 1816
79 1816
79 159
625 159
3 1 35 0 0 0 0 47 46 0 0 3
878 1810
878 1948
876 1948
2 0 9 0 0 0 0 47 0 0 149 2
869 1759
869 1304
3 1 36 0 0 8320 0 48 47 0 0 3
888 1746
887 1746
887 1759
2 0 37 0 0 4096 0 48 0 0 154 2
879 1700
879 1562
3 1 38 0 0 4224 0 49 48 0 0 2
897 1683
897 1700
1 5 39 0 0 8320 0 49 72 0 0 5
906 1638
906 1386
2126 1386
2126 275
1461 275
2 0 40 0 0 4096 0 49 0 0 153 2
888 1638
888 1588
1 0 30 0 0 0 0 50 0 0 114 2
826 1942
826 1728
0 0 30 0 0 0 0 0 0 115 0 2
826 1672
826 1732
1 0 30 0 0 8320 0 82 0 0 150 5
631 141
68 141
68 1672
826 1672
826 1329
0 1 12 0 0 0 0 0 51 151 0 2
793 1355
793 1948
3 0 14 0 0 16384 0 61 0 0 118 7
684 1324
658 1324
658 1234
44 1234
44 94
91 94
91 67
0 0 14 0 0 4224 0 0 0 0 0 3
66 67
2152 67
2152 1217
2 0 12 0 0 0 0 52 0 0 151 3
398 1388
776 1388
776 1355
3 1 41 0 0 8320 0 52 85 0 0 5
389 1339
389 1201
610 1201
610 1097
571 1097
1 1 2 0 0 4096 0 52 53 0 0 2
380 1388
380 1386
9 0 2 0 0 4096 0 85 0 0 236 2
571 1167
571 1175
1 0 2 0 0 0 0 54 0 0 162 2
571 1271
571 1272
6 11 42 0 0 4224 0 74 79 0 0 3
745 636
631 636
631 554
5 12 43 0 0 4224 0 74 79 0 0 3
745 627
613 627
613 554
13 4 44 0 0 8320 0 79 74 0 0 3
595 554
595 618
745 618
14 3 45 0 0 8320 0 79 74 0 0 3
577 554
577 609
745 609
0 14 8 0 0 4096 0 0 74 279 0 2
1053 636
809 636
0 13 7 0 0 4096 0 0 74 280 0 2
1033 627
809 627
0 12 6 0 0 4096 0 0 74 281 0 2
1013 618
809 618
0 11 5 0 0 4096 0 0 74 282 0 2
994 609
809 609
0 10 46 0 0 4096 0 0 74 283 0 2
975 600
809 600
0 9 47 0 0 4096 0 0 74 284 0 2
955 591
809 591
0 8 48 0 0 4096 0 0 74 285 0 2
935 582
809 582
0 7 49 0 0 4096 0 0 74 286 0 2
916 573
809 573
1 2 2 0 0 4224 0 75 74 0 0 2
396 600
745 600
14 3 50 0 0 4224 0 85 71 0 0 4
508 1161
508 1257
535 1257
535 1286
13 4 51 0 0 4224 0 85 71 0 0 4
517 1161
517 1262
526 1262
526 1286
12 5 52 0 0 4224 0 85 71 0 0 4
526 1161
526 1267
517 1267
517 1286
11 6 53 0 0 4224 0 85 71 0 0 4
535 1161
535 1272
508 1272
508 1286
1 0 2 0 0 0 0 91 0 0 246 3
1187 1060
1225 1060
1225 1132
1 4 54 0 0 8320 0 55 61 0 0 3
675 1357
678 1357
678 1342
3 0 9 0 0 0 0 56 0 0 149 3
736 1252
779 1252
779 1304
2 0 30 0 0 0 0 56 0 0 150 3
735 1261
774 1261
774 1329
1 0 12 0 0 0 0 56 0 0 151 3
736 1270
770 1270
770 1355
2 0 55 0 0 4096 0 61 0 0 147 3
684 1306
669 1306
669 1297
1 4 55 0 0 8320 0 61 56 0 0 4
684 1297
669 1297
669 1261
684 1261
9 1 34 0 0 12416 0 61 60 0 0 4
748 1333
766 1333
766 1278
1536 1278
10 1 9 0 0 0 0 61 57 0 0 4
748 1342
759 1342
759 1304
1536 1304
1 11 30 0 0 0 0 58 61 0 0 4
1536 1329
754 1329
754 1351
748 1351
1 12 12 0 0 0 0 59 61 0 0 4
1536 1355
754 1355
754 1360
748 1360
13 1 56 0 0 16512 0 71 69 0 0 5
562 1356
562 1610
683 1610
683 1612
1677 1612
14 1 40 0 0 24704 0 71 66 0 0 7
553 1356
553 1586
683 1586
683 1588
888 1588
888 1583
1677 1583
15 1 37 0 0 24704 0 71 65 0 0 7
544 1356
544 1560
683 1560
683 1562
879 1562
879 1560
1679 1560
16 1 22 0 0 16512 0 71 67 0 0 7
535 1356
535 1535
683 1535
683 1537
1307 1537
1307 1538
1681 1538
17 1 27 0 0 16512 0 71 68 0 0 7
526 1356
526 1509
683 1509
683 1511
1235 1511
1235 1509
1682 1509
18 1 20 0 0 0 0 71 63 0 0 7
517 1356
517 1484
684 1484
684 1486
1364 1486
1364 1485
1684 1485
19 1 18 0 0 0 0 71 64 0 0 7
508 1356
508 1458
684 1458
684 1460
1431 1460
1431 1459
1684 1459
20 1 19 0 0 0 0 71 70 0 0 5
499 1356
499 1433
684 1433
684 1435
1685 1435
21 1 33 0 0 24704 0 71 62 0 0 7
490 1356
490 1407
684 1407
684 1409
1061 1409
1061 1410
1686 1410
0 0 57 0 0 4224 0 0 0 0 0 4
684 1610
682 1610
682 1610
683 1610
1 2 2 0 0 0 0 71 71 0 0 4
571 1280
571 1272
562 1272
562 1280
0 4 58 0 0 4096 0 0 72 170 0 4
1233 316
1356 316
1356 289
1405 289
0 3 59 0 0 4096 0 0 72 169 0 4
1245 299
1343 299
1343 280
1405 280
0 2 60 0 0 4096 0 0 72 168 0 4
1255 282
1334 282
1334 271
1405 271
0 1 61 0 0 4096 0 0 72 167 0 2
1265 262
1405 262
8 8 61 0 0 8320 0 73 18 0 0 4
1228 457
1265 457
1265 262
1124 262
7 0 60 0 0 8320 0 73 0 0 270 4
1228 466
1255 466
1255 280
1134 280
6 0 59 0 0 8320 0 73 0 0 269 4
1228 475
1245 475
1245 298
1143 298
0 5 58 0 0 8320 0 0 73 268 0 4
1152 316
1236 316
1236 484
1228 484
0 0 10 0 0 0 0 0 0 0 63 2
1121 407
1126 407
0 0 10 0 0 0 0 0 0 0 63 2
1121 425
1126 425
0 0 10 0 0 0 0 0 0 0 63 2
1121 443
1126 443
2 19 62 0 0 4224 0 17 73 0 0 3
1117 452
1152 452
1152 448
4 20 63 0 0 4224 0 17 73 0 0 4
1117 434
1147 434
1147 439
1152 439
6 21 64 0 0 4224 0 17 73 0 0 4
1117 416
1142 416
1142 430
1152 430
22 8 65 0 0 12416 0 73 17 0 0 4
1152 421
1146 421
1146 398
1117 398
0 0 5 0 0 0 0 0 0 0 282 2
1057 452
994 452
0 0 6 0 0 0 0 0 0 0 281 2
1057 434
1013 434
0 0 7 0 0 0 0 0 0 0 280 2
1057 416
1033 416
12 14 66 0 0 8320 0 73 93 0 0 3
1228 421
1354 421
1354 675
11 13 67 0 0 8320 0 73 93 0 0 3
1228 430
1336 430
1336 675
10 12 68 0 0 8320 0 73 93 0 0 3
1228 439
1318 439
1318 675
9 11 69 0 0 8320 0 73 93 0 0 3
1228 448
1300 448
1300 675
8 0 49 0 0 8192 0 85 0 0 286 3
508 1097
508 935
916 935
0 7 48 0 0 4096 0 0 85 285 0 3
935 946
517 946
517 1097
6 0 47 0 0 8192 0 85 0 0 284 3
526 1097
526 961
955 961
5 0 46 0 0 8192 0 85 0 0 283 3
535 1097
535 975
975 975
2 11 70 0 0 8320 0 79 76 0 0 4
640 490
640 483
764 483
764 474
12 4 71 0 0 8320 0 76 79 0 0 4
755 474
755 480
622 480
622 490
6 13 72 0 0 8320 0 79 76 0 0 4
604 490
604 477
746 477
746 474
14 8 73 0 0 4224 0 76 79 0 0 3
737 474
586 474
586 490
5 0 8 0 0 8192 0 76 0 0 279 3
764 410
764 363
1053 363
6 0 7 0 0 8192 0 76 0 0 280 3
755 410
755 353
1033 353
7 0 6 0 0 8192 0 76 0 0 281 3
746 410
746 342
1013 342
8 0 5 0 0 8192 0 76 0 0 282 3
737 410
737 330
994 330
9 0 2 0 0 0 0 76 0 0 198 2
800 480
800 490
10 0 2 0 0 0 0 76 0 0 199 4
791 480
791 490
851 490
851 406
1 1 2 0 0 0 0 76 77 0 0 3
800 410
800 406
862 406
1 10 2 0 0 0 0 78 79 0 0 3
553 480
568 480
568 484
1 1 74 0 0 8320 0 79 2 0 0 5
649 490
649 359
263 359
263 441
218 441
1 3 75 0 0 8320 0 3 79 0 0 4
381 488
381 412
631 412
631 490
1 5 76 0 0 8320 0 4 79 0 0 4
349 487
349 397
613 397
613 490
1 7 77 0 0 8320 0 5 79 0 0 4
318 487
318 383
595 383
595 490
1 9 78 0 0 8320 0 6 79 0 0 4
285 485
285 370
577 370
577 490
0 0 5 0 0 0 0 0 0 0 282 2
858 151
994 151
0 0 6 0 0 0 0 0 0 0 281 2
858 169
1013 169
0 0 7 0 0 0 0 0 0 0 280 2
858 187
1033 187
0 0 8 0 0 0 0 0 0 0 279 2
858 205
1053 205
1 4 2 0 0 0 0 80 82 0 0 3
482 169
482 168
631 168
2 1 79 0 0 4224 0 82 81 0 0 3
631 150
598 150
598 123
0 5 5 0 0 4096 0 0 82 282 0 4
994 248
593 248
593 177
631 177
0 6 6 0 0 4096 0 0 82 281 0 4
1013 240
602 240
602 186
631 186
0 7 7 0 0 4096 0 0 82 280 0 4
1033 231
611 231
611 195
631 195
0 8 8 0 0 4096 0 0 82 279 0 4
1053 222
620 222
620 204
631 204
8 14 80 0 0 12416 0 19 82 0 0 4
797 205
794 205
794 204
695 204
0 13 13 0 0 12416 0 0 82 0 0 4
794 187
748 187
748 195
695 195
4 12 81 0 0 4224 0 19 82 0 0 4
797 169
740 169
740 186
695 186
11 2 82 0 0 12416 0 82 19 0 0 4
695 177
731 177
731 151
797 151
2 0 83 0 0 4096 0 16 0 0 263 2
1128 874
1290 874
4 0 84 0 0 4096 0 16 0 0 262 2
1128 856
1309 856
6 0 85 0 0 4224 0 16 0 0 261 2
1128 838
1327 838
8 0 86 0 0 4224 0 16 0 0 260 2
1128 820
1345 820
7 0 4 0 0 20608 0 15 0 0 80 6
812 1203
760 1203
760 1084
48 1084
48 1862
1163 1862
11 2 87 0 0 8320 0 84 15 0 0 5
664 1162
664 1186
793 1186
793 1158
818 1158
0 0 5 0 0 0 0 0 0 0 282 2
878 1212
994 1212
0 0 6 0 0 0 0 0 0 0 281 2
878 1194
1013 1194
0 0 7 0 0 0 0 0 0 0 280 2
878 1176
1033 1176
0 0 8 0 0 0 0 0 0 0 279 2
878 1158
1053 1158
12 4 88 0 0 8320 0 84 15 0 0 5
655 1162
655 1190
807 1190
807 1176
818 1176
13 6 89 0 0 8320 0 84 15 0 0 3
646 1162
646 1194
818 1194
14 0 3 0 0 8320 0 84 0 0 0 3
637 1162
637 1212
814 1212
1 0 2 0 0 0 0 83 0 0 234 4
736 1175
737 1175
737 1175
736 1175
1 0 2 0 0 0 0 84 0 0 235 4
700 1098
736 1098
736 1175
699 1175
0 9 2 0 0 0 0 0 84 236 0 3
690 1175
700 1175
700 1168
10 10 2 0 0 0 0 85 84 0 0 4
562 1167
562 1175
691 1175
691 1168
5 0 8 0 0 0 0 84 0 0 279 3
664 1098
664 1068
1053 1068
6 0 7 0 0 0 0 84 0 0 280 3
655 1098
655 1063
1033 1063
7 0 6 0 0 0 0 84 0 0 281 3
646 1098
646 1057
1013 1057
8 0 5 0 0 0 0 84 0 0 282 3
637 1098
637 1051
994 1051
11 1 90 0 0 8320 0 91 89 0 0 4
1151 1124
1151 1217
1331 1217
1331 1178
12 1 91 0 0 8320 0 91 88 0 0 4
1142 1124
1142 1210
1350 1210
1350 1178
13 1 92 0 0 8320 0 91 87 0 0 4
1133 1124
1133 1199
1370 1199
1370 1178
14 1 93 0 0 8320 0 91 86 0 0 4
1124 1124
1124 1189
1390 1189
1390 1178
9 0 2 0 0 0 0 91 0 0 246 2
1187 1130
1187 1132
10 1 2 0 0 0 0 91 90 0 0 3
1178 1130
1178 1132
1246 1132
5 0 5 0 0 0 0 91 0 0 282 3
1151 1060
1151 1036
994 1036
6 0 6 0 0 0 0 91 0 0 281 3
1142 1060
1142 1042
1013 1042
7 0 7 0 0 0 0 91 0 0 280 3
1133 1060
1133 1050
1033 1050
8 0 8 0 0 0 0 91 0 0 279 2
1124 1060
1053 1060
1 10 2 0 0 0 0 92 93 0 0 3
1393 747
1393 745
1363 745
9 0 5 0 0 0 0 16 0 0 282 2
1064 874
994 874
10 0 6 0 0 0 0 16 0 0 281 2
1064 856
1013 856
11 0 7 0 0 0 0 16 0 0 280 2
1064 838
1033 838
12 0 8 0 0 0 0 16 0 0 279 2
1064 820
1053 820
9 1 94 0 0 8320 0 93 10 0 0 4
1354 739
1354 835
1633 835
1633 955
7 1 95 0 0 8320 0 93 9 0 0 4
1336 739
1336 849
1601 849
1601 954
5 1 96 0 0 8320 0 93 8 0 0 4
1318 739
1318 864
1570 864
1570 954
3 1 97 0 0 8320 0 93 7 0 0 4
1300 739
1300 878
1537 878
1537 952
8 1 86 0 0 0 0 93 11 0 0 4
1345 739
1345 918
1386 918
1386 953
6 1 85 0 0 0 0 93 12 0 0 4
1327 739
1327 928
1354 928
1354 952
4 1 84 0 0 4224 0 93 13 0 0 4
1309 739
1309 938
1323 938
1323 952
2 1 83 0 0 8320 0 93 14 0 0 3
1291 739
1290 739
1290 950
9 0 5 0 0 0 0 18 0 0 282 2
1060 316
994 316
10 0 6 0 0 0 0 18 0 0 281 2
1060 298
1013 298
11 0 7 0 0 0 0 18 0 0 280 2
1060 280
1033 280
12 0 8 0 0 0 0 18 0 0 279 2
1060 262
1053 262
11 2 58 0 0 0 0 95 18 0 0 3
1152 234
1152 316
1124 316
12 4 59 0 0 0 0 95 18 0 0 3
1143 234
1143 298
1124 298
13 6 60 0 0 0 0 95 18 0 0 3
1134 234
1134 280
1124 280
14 0 61 0 0 0 0 95 0 0 167 3
1125 234
1128 234
1128 262
1 0 2 0 0 0 0 95 0 0 274 3
1188 170
1220 170
1220 243
9 0 2 0 0 0 0 95 0 0 274 2
1188 240
1188 243
10 1 2 0 0 0 0 95 94 0 0 3
1179 240
1179 243
1247 243
5 0 5 0 0 0 0 95 0 0 282 3
1152 170
1152 146
994 146
6 0 6 0 0 0 0 95 0 0 281 3
1143 170
1143 152
1013 152
7 0 7 0 0 0 0 95 0 0 280 3
1134 170
1134 160
1033 160
8 0 8 0 0 0 0 95 0 0 279 2
1125 170
1053 170
1 1 8 0 0 4224 0 107 100 0 0 2
1053 112
1053 1225
1 1 7 0 0 4224 0 106 101 0 0 2
1033 112
1033 1225
1 1 6 0 0 4224 0 105 102 0 0 2
1013 112
1013 1225
1 1 5 0 0 4224 0 104 103 0 0 2
994 112
994 1225
1 1 46 0 0 4224 0 108 99 0 0 2
975 112
975 1225
1 1 47 0 0 4224 0 109 98 0 0 2
955 112
955 1225
1 1 48 0 0 4224 0 110 97 0 0 2
935 112
935 1225
1 1 49 0 0 4224 0 111 96 0 0 2
916 112
916 1225
56
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
190 446 288 469
202 456 275 471
9 SM(MAR=1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
704 1588 755 1611
717 1598 741 1613
3 HLT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
708 1565 751 1588
721 1575 737 1590
2 JZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1537 757 1560
720 1547 744 1562
3 JMP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1514 757 1537
720 1524 744 1539
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
707 1488 758 1511
720 1498 744 1513
3 MOV
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1460 757 1483
720 1470 744 1485
3 AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
706 1436 757 1459
719 1446 743 1461
3 SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
708 1409 757 1432
720 1419 744 1434
3 ADD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
709 1382 758 1405
721 1392 745 1407
3 LDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 1331 833 1354
803 1341 819 1356
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 1304 829 1327
800 1314 816 1329
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
789 1280 832 1303
802 1290 818 1305
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 1252 833 1275
803 1262 819 1277
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
704 96 739 118
713 103 729 119
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
809 364 852 386
818 371 842 387
3 MAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
420 418 527 440
429 425 517 441
11 INPUT & MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
755 652 798 674
764 660 788 676
3 RAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
654 986 689 1008
663 994 679 1010
2 IR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1275 201 1304 223
1285 208 1293 224
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1373 426 1416 448
1382 434 1406 450
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1409 699 1452 721
1418 706 1442 722
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1163 919 1190 941
1172 926 1180 942
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1504 913 1531 935
1513 920 1521 936
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1229 1051 1304 1073
1238 1058 1294 1074
7 OUT REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1418 1148 1493 1170
1427 1155 1483 1171
7 DISPLAY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
79 30 123 54
90 39 111 55
3 clk
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
778 73 815 97
789 81 803 97
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
758 1963 795 1987
769 1971 783 1987
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
811 1965 848 1989
822 1974 836 1990
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
493 113 530 137
504 122 518 138
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
861 1974 898 1998
872 1983 886 1999
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
126 167 157 191
134 176 148 192
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
931 2001 964 2025
940 2010 954 2026
2 Lm
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1030 2007 1063 2031
1039 2016 1053 2032
2 Cs
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
797 289 834 313
808 298 822 314
2 Lm
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
335 538 368 562
344 547 358 563
2 Cs
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1101 2004 1134 2028
1110 2012 1124 2028
2 Li
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
290 988 327 1012
301 997 315 1013
2 Li
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1147 1994 1184 2018
1158 2003 1172 2019
2 Ei
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1216 2000 1253 2024
1227 2009 1241 2025
2 La
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1290 126 1327 150
1301 135 1315 151
2 La
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1287 2021 1324 2045
1298 2030 1312 2046
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1971 330 2002 354
1979 339 1993 355
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1968 386 2005 410
1979 393 1993 409
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1434 2049 1467 2073
1443 2058 1457 2074
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1348 2042 1385 2066
1359 2050 1373 2066
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1423 2067 1460 2091
1434 2076 1448 2092
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1483 2052 1516 2076
1492 2060 1506 2076
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1536 1654 1569 1678
1545 1662 1559 1678
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1564 1676 1588 1700
1572 1685 1579 1701
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1570 1705 1614 1729
1581 1714 1602 1730
3 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1606 2118 1643 2142
1617 2127 1631 2143
2 Eb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1699 2127 1736 2151
1710 2136 1724 2152
2 Lo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1809 813 1846 837
1820 822 1834 838
2 Eb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1752 981 1789 1005
1763 990 1777 1006
2 Lo
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
