CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
48
13 Logic Switch~
5 609 105 0 1 11
0 3
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V33
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4244 0 0
2
42919.8 0
0
13 Logic Switch~
5 635 114 0 1 11
0 2
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V37
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5225 0 0
2
42919.8 0
0
13 Logic Switch~
5 777 96 0 1 11
0 4
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V35
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
768 0 0
2
42919.8 0
0
13 Logic Switch~
5 601 87 0 1 11
0 5
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V34
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5735 0 0
2
42919.8 0
0
13 Logic Switch~
5 22 562 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V32
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5881 0 0
2
42919.8 7
0
13 Logic Switch~
5 27 588 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V31
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3275 0 0
2
42919.8 6
0
13 Logic Switch~
5 29 603 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V30
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4203 0 0
2
42919.8 5
0
13 Logic Switch~
5 30 624 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V29
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3440 0 0
2
42919.8 4
0
13 Logic Switch~
5 26 641 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V28
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9102 0 0
2
42919.8 3
0
13 Logic Switch~
5 25 654 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V27
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5586 0 0
2
42919.8 2
0
13 Logic Switch~
5 26 667 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V26
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
525 0 0
2
42919.8 1
0
13 Logic Switch~
5 26 691 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V25
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6206 0 0
2
42919.8 0
0
13 Logic Switch~
5 22 391 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V24
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3418 0 0
2
42919.8 7
0
13 Logic Switch~
5 27 417 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V23
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9312 0 0
2
42919.8 6
0
13 Logic Switch~
5 29 432 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V22
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7419 0 0
2
42919.8 5
0
13 Logic Switch~
5 30 453 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V21
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
472 0 0
2
42919.8 4
0
13 Logic Switch~
5 26 470 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4714 0 0
2
42919.8 3
0
13 Logic Switch~
5 25 483 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9386 0 0
2
42919.8 2
0
13 Logic Switch~
5 26 496 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7610 0 0
2
42919.8 1
0
13 Logic Switch~
5 26 520 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3482 0 0
2
42919.8 0
0
13 Logic Switch~
5 19 213 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3608 0 0
2
42919.8 7
0
13 Logic Switch~
5 24 239 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6397 0 0
2
42919.8 6
0
13 Logic Switch~
5 26 254 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3967 0 0
2
42919.8 5
0
13 Logic Switch~
5 27 275 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8621 0 0
2
42919.8 4
0
13 Logic Switch~
5 23 292 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
42919.8 3
0
13 Logic Switch~
5 22 305 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7385 0 0
2
42919.8 2
0
13 Logic Switch~
5 23 318 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6519 0 0
2
42919.8 1
0
13 Logic Switch~
5 23 342 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
552 0 0
2
42919.8 0
0
13 Logic Switch~
5 28 149 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5551 0 0
2
42919.8 0
0
13 Logic Switch~
5 28 125 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8715 0 0
2
42919.8 0
0
13 Logic Switch~
5 27 112 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9763 0 0
2
42919.8 0
0
13 Logic Switch~
5 28 99 0 1 11
0 41
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8443 0 0
2
42919.8 0
0
13 Logic Switch~
5 32 82 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3719 0 0
2
42919.8 0
0
13 Logic Switch~
5 31 61 0 1 11
0 43
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8671 0 0
2
42919.8 0
0
13 Logic Switch~
5 29 46 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
42919.8 0
0
13 Logic Switch~
5 24 20 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
49 0 0
2
42919.8 0
0
14 Logic Display~
6 601 689 0 1 2
10 6
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L9
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6536 0 0
2
42919.8 0
0
14 Logic Display~
6 731 680 0 1 2
10 7
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3931 0 0
2
42919.8 0
0
14 Logic Display~
6 735 509 0 1 2
10 8
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4390 0 0
2
42919.8 0
0
14 Logic Display~
6 608 518 0 1 2
10 9
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3242 0 0
2
42919.8 0
0
14 Logic Display~
6 603 340 0 1 2
10 10
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6760 0 0
2
42919.8 0
0
14 Logic Display~
6 750 331 0 1 2
10 11
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5760 0 0
2
42919.8 0
0
14 Logic Display~
6 617 147 0 1 2
10 12
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3781 0 0
2
42919.8 0
0
14 Logic Display~
6 723 138 0 1 2
10 13
0
0 0 53856 602
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8545 0 0
2
42919.8 0
0
7 74LS151
20 296 656 0 14 29
0 21 20 19 18 17 16 15 14 5
4 3 2 7 6
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
9739 0 0
2
42919.8 8
0
7 74LS151
20 296 485 0 14 29
0 29 28 27 26 25 24 23 22 5
4 3 2 8 9
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
388 0 0
2
42919.8 8
0
7 74LS151
20 293 307 0 14 29
0 37 36 35 34 33 32 31 30 5
4 3 2 11 10
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
4595 0 0
2
42919.8 8
0
7 74LS151
20 298 114 0 14 29
0 45 44 43 42 41 40 39 38 5
4 3 2 13 12
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
3173 0 0
2
42919.8 0
0
100
0 0 2 0 0 4096 0 0 0 10 89 2
477 310
477 114
0 0 3 0 0 4096 0 0 0 11 90 2
504 302
504 105
0 0 4 0 0 4096 0 0 0 12 91 2
534 292
534 96
0 0 5 0 0 4096 0 0 0 13 92 2
559 280
559 87
1 0 3 0 0 0 0 1 0 0 90 2
597 105
597 105
12 12 2 0 0 0 0 46 45 0 0 4
328 485
477 485
477 656
328 656
11 11 3 0 0 0 0 46 45 0 0 4
328 476
504 476
504 647
328 647
10 10 4 0 0 4096 0 46 45 0 0 4
328 467
534 467
534 638
328 638
9 9 5 0 0 4096 0 46 45 0 0 4
334 458
561 458
561 629
334 629
12 0 2 0 0 0 0 47 0 0 6 3
325 307
477 307
477 489
11 0 3 0 0 0 0 47 0 0 7 3
325 298
504 298
504 476
10 0 4 0 0 4096 0 47 0 0 8 3
325 289
534 289
534 470
9 0 5 0 0 4096 0 47 0 0 9 3
331 280
560 280
560 458
1 0 6 0 0 0 0 37 0 0 33 2
586 692
586 692
1 0 7 0 0 0 0 38 0 0 34 2
716 683
716 683
1 0 8 0 0 0 0 39 0 0 52 2
720 512
720 512
1 0 9 0 0 0 0 40 0 0 51 2
593 521
593 521
1 0 10 0 0 0 0 41 0 0 69 2
588 343
588 343
1 0 11 0 0 0 0 42 0 0 70 2
735 334
735 334
1 0 12 0 0 0 0 43 0 0 87 2
602 150
602 150
1 0 13 0 0 0 0 44 0 0 88 2
708 141
708 141
1 0 2 0 0 0 0 2 0 0 89 2
623 114
623 114
1 0 4 0 0 0 0 3 0 0 91 2
765 96
765 96
1 0 5 0 0 0 0 4 0 0 92 2
589 87
589 87
1 0 14 0 0 4096 0 12 0 0 35 2
38 691
38 692
1 0 15 0 0 0 0 11 0 0 36 2
38 667
38 667
1 0 16 0 0 0 0 10 0 0 37 2
37 654
37 654
1 0 17 0 0 0 0 9 0 0 38 2
38 641
38 641
1 0 18 0 0 0 0 8 0 0 39 2
42 624
42 624
1 0 19 0 0 0 0 7 0 0 40 2
41 603
41 603
1 0 20 0 0 0 0 6 0 0 41 2
39 588
39 588
1 0 21 0 0 0 0 5 0 0 42 2
34 562
34 562
14 0 6 0 0 4224 0 45 0 0 0 2
334 692
604 692
13 0 7 0 0 4224 0 45 0 0 0 2
328 683
733 683
8 0 14 0 0 4224 0 45 0 0 0 2
264 692
22 692
7 0 15 0 0 4224 0 45 0 0 0 4
264 683
72 683
72 667
22 667
6 0 16 0 0 4224 0 45 0 0 0 4
264 674
84 674
84 654
23 654
5 0 17 0 0 4224 0 45 0 0 0 4
264 665
94 665
94 641
22 641
4 0 18 0 0 4224 0 45 0 0 0 4
264 656
108 656
108 624
22 624
3 0 19 0 0 4224 0 45 0 0 0 4
264 647
121 647
121 603
19 603
2 0 20 0 0 4224 0 45 0 0 0 4
264 638
135 638
135 588
22 588
1 0 21 0 0 12416 0 45 0 0 0 4
264 629
150 629
150 562
27 562
1 0 22 0 0 4096 0 20 0 0 53 2
38 520
38 521
1 0 23 0 0 0 0 19 0 0 54 2
38 496
38 496
1 0 24 0 0 0 0 18 0 0 55 2
37 483
37 483
1 0 25 0 0 0 0 17 0 0 56 2
38 470
38 470
1 0 26 0 0 0 0 16 0 0 57 2
42 453
42 453
1 0 27 0 0 0 0 15 0 0 58 2
41 432
41 432
1 0 28 0 0 0 0 14 0 0 59 2
39 417
39 417
1 0 29 0 0 0 0 13 0 0 60 2
34 391
34 391
14 0 9 0 0 4224 0 46 0 0 0 2
334 521
604 521
13 0 8 0 0 4224 0 46 0 0 0 2
328 512
735 512
8 0 22 0 0 4224 0 46 0 0 0 2
264 521
22 521
7 0 23 0 0 4224 0 46 0 0 0 4
264 512
72 512
72 496
22 496
6 0 24 0 0 4224 0 46 0 0 0 4
264 503
84 503
84 483
23 483
5 0 25 0 0 4224 0 46 0 0 0 4
264 494
94 494
94 470
22 470
4 0 26 0 0 4224 0 46 0 0 0 4
264 485
108 485
108 453
22 453
3 0 27 0 0 4224 0 46 0 0 0 4
264 476
121 476
121 432
19 432
2 0 28 0 0 4224 0 46 0 0 0 4
264 467
135 467
135 417
22 417
1 0 29 0 0 12416 0 46 0 0 0 4
264 458
150 458
150 391
27 391
1 0 30 0 0 4096 0 28 0 0 71 2
35 342
35 343
1 0 31 0 0 0 0 27 0 0 72 2
35 318
35 318
1 0 32 0 0 0 0 26 0 0 73 2
34 305
34 305
1 0 33 0 0 0 0 25 0 0 74 2
35 292
35 292
1 0 34 0 0 0 0 24 0 0 75 2
39 275
39 275
1 0 35 0 0 0 0 23 0 0 76 2
38 254
38 254
1 0 36 0 0 0 0 22 0 0 77 2
36 239
36 239
1 0 37 0 0 0 0 21 0 0 78 2
31 213
31 213
14 0 10 0 0 4224 0 47 0 0 0 3
331 343
598 343
598 345
13 0 11 0 0 4224 0 47 0 0 0 2
325 334
741 334
8 0 30 0 0 4224 0 47 0 0 0 2
261 343
19 343
7 0 31 0 0 4224 0 47 0 0 0 4
261 334
69 334
69 318
19 318
6 0 32 0 0 4224 0 47 0 0 0 4
261 325
81 325
81 305
20 305
5 0 33 0 0 4224 0 47 0 0 0 4
261 316
91 316
91 292
19 292
4 0 34 0 0 4224 0 47 0 0 0 4
261 307
105 307
105 275
19 275
3 0 35 0 0 4224 0 47 0 0 0 4
261 298
118 298
118 254
16 254
2 0 36 0 0 4224 0 47 0 0 0 4
261 289
132 289
132 239
19 239
1 0 37 0 0 12416 0 47 0 0 0 4
261 280
147 280
147 213
24 213
1 0 38 0 0 4096 0 29 0 0 93 2
40 149
40 150
1 0 39 0 0 0 0 30 0 0 94 2
40 125
40 125
1 0 40 0 0 0 0 31 0 0 95 2
39 112
39 112
1 0 41 0 0 0 0 32 0 0 96 2
40 99
40 99
1 0 42 0 0 0 0 33 0 0 97 2
44 82
44 82
1 0 43 0 0 0 0 34 0 0 98 2
43 61
43 61
1 0 44 0 0 0 0 35 0 0 99 2
41 46
41 46
1 0 45 0 0 0 0 36 0 0 100 2
36 20
36 20
14 0 12 0 0 4224 0 48 0 0 0 2
336 150
606 150
13 0 13 0 0 4224 0 48 0 0 0 2
330 141
713 141
12 0 2 0 0 4224 0 48 0 0 0 2
330 114
638 114
11 0 3 0 0 4224 0 48 0 0 0 2
330 105
606 105
10 0 4 0 0 4224 0 48 0 0 0 2
330 96
781 96
9 0 5 0 0 4224 0 48 0 0 0 2
336 87
605 87
8 0 38 0 0 4224 0 48 0 0 0 2
266 150
24 150
7 0 39 0 0 4224 0 48 0 0 0 4
266 141
74 141
74 125
24 125
6 0 40 0 0 4224 0 48 0 0 0 4
266 132
86 132
86 112
25 112
5 0 41 0 0 4224 0 48 0 0 0 4
266 123
96 123
96 99
24 99
4 0 42 0 0 4224 0 48 0 0 0 4
266 114
110 114
110 82
24 82
3 0 43 0 0 4224 0 48 0 0 0 4
266 105
123 105
123 61
21 61
2 0 44 0 0 4224 0 48 0 0 0 4
266 96
137 96
137 46
24 46
1 0 45 0 0 12416 0 48 0 0 0 4
266 87
152 87
152 20
29 20
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
