CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
27
7 Ground~
168 938 102 0 1 3
0 0
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
42655.5 0
0
7 74LS173
129 462 112 0 1 29
0 0
0
0 0 4832 0
7 74LS173
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
391 0 0
2
42655.5 25
0
7 74LS173
129 603 104 0 1 29
0 0
0
0 0 4832 0
7 74LS173
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
3124 0 0
2
42655.5 24
0
6 Diode~
219 399 277 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
3421 0 0
2
42655.5 23
0
6 Diode~
219 454 275 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D2
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
8157 0 0
2
42655.5 22
0
6 Diode~
219 511 274 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D3
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
5572 0 0
2
42655.5 21
0
6 Diode~
219 568 274 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D4
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
8901 0 0
2
42655.5 20
0
6 Diode~
219 827 271 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D5
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
7361 0 0
2
42655.5 19
0
6 Diode~
219 770 271 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D6
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
4747 0 0
2
42655.5 18
0
6 Diode~
219 713 272 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D7
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
972 0 0
2
42655.5 17
0
6 Diode~
219 658 274 0 1 5
0 0
0
0 0 832 270
5 DIODE
11 0 46 8
2 D8
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
3472 0 0
2
42655.5 16
0
9 Resistor~
219 400 223 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9998 0 0
2
42655.5 15
0
9 Resistor~
219 453 228 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3536 0 0
2
42655.5 14
0
9 Resistor~
219 510 227 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4597 0 0
2
42655.5 13
0
9 Resistor~
219 568 232 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3835 0 0
2
42655.5 12
0
9 Resistor~
219 822 221 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3670 0 0
2
42655.5 11
0
9 Resistor~
219 764 216 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5616 0 0
2
42655.5 10
0
9 Resistor~
219 707 217 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9323 0 0
2
42655.5 9
0
9 Resistor~
219 654 212 0 1 5
0 0
0
0 0 864 782
2 1k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
317 0 0
2
42655.5 8
0
7 Ground~
168 399 313 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3108 0 0
2
42655.5 7
0
7 Ground~
168 452 315 0 1 3
0 0
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4299 0 0
2
42655.5 6
0
7 Ground~
168 511 317 0 1 3
0 0
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9672 0 0
2
42655.5 5
0
7 Ground~
168 569 315 0 1 3
0 0
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7876 0 0
2
42655.5 4
0
7 Ground~
168 832 314 0 1 3
0 0
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6369 0 0
2
42655.5 3
0
7 Ground~
168 774 316 0 1 3
0 0
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9172 0 0
2
42655.5 2
0
7 Ground~
168 715 314 0 1 3
0 0
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7100 0 0
2
42655.5 1
0
7 Ground~
168 662 312 0 1 3
0 0
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3820 0 0
2
42655.5 0
0
52
4 0 0 0 0 0 0 3 0 0 2 3
571 104
560 104
560 258
4 0 0 0 0 0 0 2 0 0 0 9
430 112
420 112
420 258
758 258
758 284
937 284
937 258
951 258
951 266
0 0 0 0 0 0 0 0 0 7 4 3
565 90
645 90
645 47
0 1 0 0 0 0 0 0 1 5 0 5
424 99
415 99
415 47
938 47
938 96
3 2 0 0 0 0 0 2 2 0 0 2
424 103
424 94
3 2 0 0 0 0 0 2 2 0 0 2
424 103
424 94
3 2 0 0 0 0 0 3 3 0 0 2
565 95
565 86
1 0 0 0 0 0 0 2 0 0 9 4
430 85
420 85
420 58
561 58
1 0 0 0 0 0 0 3 0 0 10 3
571 77
561 77
561 57
0 0 0 0 0 0 0 0 0 13 11 5
500 89
561 89
561 57
833 57
833 86
10 0 0 0 0 0 0 3 0 0 0 3
641 86
885 86
885 124
10 9 0 0 0 0 0 3 3 0 0 2
641 86
641 77
10 9 0 0 0 0 0 2 2 0 0 2
500 94
500 85
5 0 0 0 0 0 0 3 0 0 24 3
571 113
571 161
309 161
6 0 0 0 0 0 0 3 0 0 28 6
571 122
521 122
521 39
324 39
324 109
282 109
7 0 0 0 0 0 0 3 0 0 23 6
571 131
529 131
529 56
331 56
331 213
256 213
8 0 0 0 0 0 0 3 0 0 27 6
571 140
543 140
543 50
351 50
351 227
229 227
5 0 0 0 0 0 0 2 0 0 22 4
430 121
316 121
316 251
200 251
6 0 0 0 0 0 0 2 0 0 26 4
430 130
321 130
321 263
171 263
7 0 0 0 0 0 0 2 0 0 21 4
430 139
340 139
340 284
142 284
0 0 0 0 0 0 0 0 0 0 0 2
142 293
142 56
0 0 0 0 0 0 0 0 0 0 0 2
200 293
200 69
0 0 0 0 0 0 0 0 0 0 0 2
256 290
256 60
0 0 0 0 0 0 0 0 0 0 0 2
309 291
309 61
8 0 0 0 0 0 0 2 0 0 0 6
430 148
370 148
370 301
115 301
115 45
117 45
0 0 0 0 0 0 0 0 0 0 0 2
171 55
171 293
0 0 0 0 0 0 0 0 0 0 0 2
229 57
229 290
0 0 0 0 0 0 0 0 0 0 0 2
282 60
282 291
1 2 0 0 0 0 0 24 8 0 0 4
832 308
832 289
827 289
827 281
1 2 0 0 0 0 0 25 9 0 0 4
774 310
774 289
770 289
770 281
1 2 0 0 0 0 0 26 10 0 0 4
715 308
715 290
713 290
713 282
1 2 0 0 0 0 0 27 11 0 0 4
662 306
662 292
658 292
658 284
1 2 0 0 0 0 0 23 7 0 0 4
569 309
569 292
568 292
568 284
1 2 0 0 0 0 0 22 6 0 0 2
511 311
511 284
1 2 0 0 0 0 0 21 5 0 0 4
452 309
452 293
454 293
454 285
1 2 0 0 0 0 0 20 4 0 0 2
399 307
399 287
2 1 0 0 0 0 0 12 4 0 0 4
400 241
400 259
399 259
399 267
14 1 0 0 0 0 0 2 12 0 0 5
494 148
463 148
463 197
400 197
400 205
2 1 0 0 0 0 0 13 5 0 0 4
453 246
453 257
454 257
454 265
13 1 0 0 0 0 0 2 13 0 0 5
494 139
458 139
458 202
453 202
453 210
2 1 0 0 0 0 0 14 6 0 0 4
510 245
510 256
511 256
511 264
12 1 0 0 0 0 0 2 14 0 0 3
494 130
510 130
510 209
2 1 0 0 0 0 0 15 7 0 0 2
568 250
568 264
11 1 0 0 0 0 0 2 15 0 0 5
494 121
538 121
538 200
568 200
568 214
2 1 0 0 0 0 0 19 11 0 0 4
654 230
654 256
658 256
658 264
14 1 0 0 0 0 0 3 19 0 0 3
635 140
654 140
654 194
2 1 0 0 0 0 0 18 10 0 0 4
707 235
707 254
713 254
713 262
13 1 0 0 0 0 0 3 18 0 0 3
635 131
707 131
707 199
2 1 0 0 0 0 0 17 9 0 0 4
764 234
764 253
770 253
770 261
12 1 0 0 0 0 0 3 17 0 0 3
635 122
764 122
764 198
2 1 0 0 0 0 0 16 8 0 0 4
822 239
822 253
827 253
827 261
11 1 0 0 0 0 0 3 16 0 0 3
635 113
822 113
822 203
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
870 136 911 157
878 143 902 158
3 Lo'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
947 278 988 299
955 285 979 300
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
111 19 306 63
116 23 300 55
23 I7 I6 I5 I4 I3 I2 I1 I0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
602 24 743 48
612 32 732 48
15 OUTPUT REGISTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
