CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
69
13 Logic Switch~
5 907 33 0 10 11
0 62 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8324 0 0
2
42920 0
0
13 Logic Switch~
5 408 35 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9550 0 0
2
42920 0
0
13 Logic Switch~
5 375 34 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6380 0 0
2
42920 0
0
13 Logic Switch~
5 337 35 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7942 0 0
2
42920 0
0
13 Logic Switch~
5 302 35 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
789 0 0
2
42920 0
0
13 Logic Switch~
5 266 35 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9884 0 0
2
42920 0
0
13 Logic Switch~
5 232 34 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6253 0 0
2
42920 0
0
13 Logic Switch~
5 25 35 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7409 0 0
2
42920 0
0
13 Logic Switch~
5 91 35 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3540 0 0
2
42920 0
0
13 Logic Switch~
5 146 34 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
10 -30 24 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3103 0 0
2
42920 0
0
9 Inverter~
13 629 1424 0 2 22
0 3 6
0
0 0 624 692
6 74LS04
-21 -19 21 -11
4 U25E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 25 0
1 U
3548 0 0
2
42920.7 0
0
9 Inverter~
13 632 1062 0 2 22
0 4 7
0
0 0 624 692
6 74LS04
-21 -19 21 -11
4 U25D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 25 0
1 U
9961 0 0
2
42920.7 0
0
9 Inverter~
13 643 724 0 2 22
0 5 8
0
0 0 624 692
6 74LS04
-21 -19 21 -11
4 U25C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 25 0
1 U
8521 0 0
2
42920.7 0
0
9 Inverter~
13 652 384 0 2 22
0 2 9
0
0 0 624 692
6 74LS04
-21 -19 21 -11
4 U25A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 25 0
1 U
5296 0 0
2
42920.7 0
0
8 4-In OR~
219 660 622 0 5 22
0 30 31 32 33 54
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U24A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 24 0
1 U
5398 0 0
2
42920.6 0
0
14 Logic Display~
6 1107 175 0 1 2
10 66
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7935 0 0
2
42920 0
0
14 Logic Display~
6 1142 176 0 1 2
10 64
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
356 0 0
2
42920 0
0
14 Logic Display~
6 1189 175 0 1 2
10 65
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4629 0 0
2
42920 0
0
14 Logic Display~
6 1227 173 0 1 2
10 63
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
2
42920 0
0
5 4071~
219 802 1174 0 3 22
0 51 50 61
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U23D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 23 0
1 U
5713 0 0
2
42920 0
0
5 4071~
219 796 870 0 3 22
0 53 52 60
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U23C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 23 0
1 U
6618 0 0
2
42920 0
0
5 4071~
219 789 520 0 3 22
0 55 54 59
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U23B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 23 0
1 U
3714 0 0
2
42920 0
0
5 4071~
219 788 186 0 3 22
0 57 56 58
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U23A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 23 0
1 U
9116 0 0
2
42920 0
0
9 2-In AND~
219 976 189 0 3 22
0 58 62 66
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U22A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
7960 0 0
2
42920 4
0
9 2-In AND~
219 993 516 0 3 22
0 59 62 64
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U22B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
3886 0 0
2
42920 3
0
9 2-In AND~
219 985 854 0 3 22
0 60 62 65
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U22C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 22 0
1 U
3299 0 0
2
42920 2
0
9 2-In AND~
219 1008 1192 0 3 22
0 61 62 63
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U22D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 22 0
1 U
9107 0 0
2
42920 1
0
8 4-In OR~
219 669 1300 0 5 22
0 47 46 48 49 50
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U21B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 21 0
1 U
6556 0 0
2
42920 0
0
8 4-In OR~
219 669 1140 0 5 22
0 42 43 44 45 51
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U21A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 21 0
1 U
3205 0 0
2
42920 0
0
8 4-In OR~
219 667 961 0 5 22
0 34 36 38 40 52
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U20B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 20 0
1 U
7255 0 0
2
42920 0
0
8 4-In OR~
219 666 804 0 5 22
0 41 39 37 35 53
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U20A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 20 0
1 U
8613 0 0
2
42920 0
0
8 4-In OR~
219 665 457 0 5 22
0 29 28 27 26 55
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U19A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 19 0
1 U
7832 0 0
2
42920 0
0
8 4-In OR~
219 661 290 0 5 22
0 21 20 19 18 56
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 18 0
1 U
8937 0 0
2
42920 0
0
8 4-In OR~
219 674 119 0 5 22
0 25 24 23 22 57
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 18 0
1 U
556 0 0
2
42920 0
0
5 4082~
219 490 694 0 5 22
0 5 14 10 11 33
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
6981 0 0
2
42920 23
0
5 4082~
219 490 653 0 5 22
0 8 14 10 12 32
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
8701 0 0
2
42920 22
0
5 4082~
219 490 612 0 5 22
0 2 14 13 11 31
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
5540 0 0
2
42920 21
0
5 4082~
219 490 572 0 5 22
0 4 14 13 12 30
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
8365 0 0
2
42920 20
0
5 4082~
219 491 531 0 5 22
0 2 15 10 11 26
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
5209 0 0
2
42920 19
0
5 4082~
219 491 491 0 5 22
0 4 15 10 12 27
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
3297 0 0
2
42920 18
0
5 4082~
219 492 451 0 5 22
0 17 15 13 67 28
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 9 0
1 U
9904 0 0
2
42920 17
0
5 4082~
219 493 410 0 5 22
0 16 15 13 12 29
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
6918 0 0
2
42920 16
0
5 4082~
219 487 1037 0 5 22
0 4 14 10 11 40
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
7751 0 0
2
42920 15
0
5 4082~
219 487 996 0 5 22
0 7 14 10 12 38
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
9907 0 0
2
42920 14
0
5 4082~
219 487 955 0 5 22
0 5 14 13 11 36
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U11A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 11 0
1 U
6628 0 0
2
42920 13
0
5 4082~
219 487 915 0 5 22
0 3 14 13 12 34
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U11B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 11 0
1 U
4914 0 0
2
42920 12
0
5 4082~
219 488 874 0 5 22
0 5 15 10 11 35
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U12A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
635 0 0
2
42920 11
0
5 4082~
219 488 834 0 5 22
0 3 15 10 12 37
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U12B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 12 0
1 U
3606 0 0
2
42920 10
0
5 4082~
219 489 794 0 5 22
0 17 15 13 11 39
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U13A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
8769 0 0
2
42920 9
0
5 4082~
219 490 753 0 5 22
0 16 15 13 12 41
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U13B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
3887 0 0
2
42920 8
0
5 4082~
219 485 1385 0 5 22
0 3 14 10 11 49
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
4266 0 0
2
42920 7
0
5 4082~
219 485 1344 0 5 22
0 6 14 10 12 48
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
3389 0 0
2
42920 6
0
5 4082~
219 485 1303 0 5 22
0 4 14 13 11 46
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 15 0
1 U
8108 0 0
2
42920 5
0
5 4082~
219 485 1263 0 5 22
0 17 14 13 12 47
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 15 0
1 U
3301 0 0
2
42920 4
0
5 4082~
219 486 1222 0 5 22
0 4 15 10 11 45
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
3739 0 0
2
42920 3
0
5 4082~
219 486 1182 0 5 22
0 2 15 10 12 44
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 16 0
1 U
4610 0 0
2
42920 2
0
5 4082~
219 487 1142 0 5 22
0 17 15 13 11 43
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U17A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 17 0
1 U
7104 0 0
2
42920 1
0
5 4082~
219 488 1101 0 5 22
0 16 15 13 12 42
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U17B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 17 0
1 U
5233 0 0
2
42920 0
0
5 4082~
219 493 359 0 5 22
0 2 14 10 11 18
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
345 0 0
2
42920 7
0
5 4082~
219 493 318 0 5 22
0 9 14 10 12 19
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
4311 0 0
2
42920 6
0
5 4082~
219 493 277 0 5 22
0 17 14 13 11 20
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
3959 0 0
2
42920 5
0
5 4082~
219 493 237 0 5 22
0 5 14 13 12 21
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
9550 0 0
2
42920 4
0
5 4082~
219 494 196 0 5 22
0 3 10 11 15 22
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
4183 0 0
2
42920 3
0
5 4082~
219 494 156 0 5 22
0 5 15 10 12 23
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
7662 0 0
2
42920 2
0
5 4082~
219 495 116 0 5 22
0 17 15 13 11 24
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
6373 0 0
2
42920 1
0
5 4082~
219 496 75 0 5 22
0 16 15 13 12 25
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
76 0 0
2
42920 0
0
9 Inverter~
13 39 48 0 2 22
0 15 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
4168 0 0
2
42920 0
0
9 Inverter~
13 105 49 0 2 22
0 13 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
9490 0 0
2
42920 0
0
9 Inverter~
13 162 51 0 2 22
0 12 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
3202 0 0
2
42920 0
0
211
0 0 2 0 0 12416 0 0 0 64 203 6
418 1169
418 1499
197 1499
197 339
318 339
318 346
0 0 3 0 0 4096 0 0 0 87 200 2
380 821
380 1372
0 0 4 0 0 4096 0 0 0 107 201 2
366 478
366 1024
0 0 5 0 0 4096 0 0 0 127 202 2
390 143
390 681
0 0 3 0 0 12288 0 0 0 200 126 6
429 1372
429 1475
210 1475
210 178
287 178
287 183
0 0 4 0 0 0 0 0 0 201 63 2
389 1024
389 1209
0 0 5 0 0 0 0 0 0 202 86 2
400 681
400 861
0 0 2 0 0 0 0 0 0 203 104 2
426 346
426 518
0 0 3 0 0 0 0 0 0 85 200 2
398 902
398 1372
0 0 4 0 0 0 0 0 0 101 201 2
425 559
425 1024
0 0 5 0 0 0 0 0 0 125 202 2
432 224
432 681
0 0 2 0 0 0 0 0 0 100 203 2
453 599
453 346
0 0 5 0 0 0 0 0 0 84 202 2
453 942
453 681
0 0 4 0 0 0 0 0 0 62 201 2
441 1290
441 1024
2 0 6 0 0 8320 0 11 0 0 61 4
650 1424
650 1447
269 1447
269 1331
0 1 3 0 0 0 0 0 11 200 0 3
439 1372
439 1424
614 1424
2 0 7 0 0 8320 0 12 0 0 83 4
653 1062
653 1072
261 1072
261 983
0 1 4 0 0 0 0 0 12 201 0 3
451 1024
451 1062
617 1062
2 0 8 0 0 8320 0 13 0 0 99 4
664 724
664 735
289 735
289 640
0 1 5 0 0 0 0 0 13 202 0 3
439 681
439 724
628 724
2 0 9 0 0 8320 0 14 0 0 118 4
673 384
673 392
243 392
243 305
0 1 2 0 0 0 0 0 14 203 0 3
442 346
442 384
637 384
3 0 10 0 0 4096 0 59 0 0 41 2
469 364
126 364
3 0 10 0 0 0 0 60 0 0 41 2
469 323
126 323
2 0 10 0 0 4096 0 63 0 0 41 2
470 192
126 192
3 0 10 0 0 0 0 64 0 0 41 2
470 161
126 161
4 0 11 0 0 4096 0 35 0 0 204 2
466 708
183 708
3 0 10 0 0 0 0 35 0 0 41 2
466 699
126 699
3 0 10 0 0 0 0 36 0 0 41 2
466 658
126 658
3 0 10 0 0 0 0 39 0 0 41 2
467 536
126 536
3 0 10 0 0 0 0 40 0 0 41 2
467 496
126 496
3 0 10 0 0 0 0 47 0 0 41 2
464 879
126 879
3 0 10 0 0 0 0 48 0 0 41 2
464 839
126 839
3 0 10 0 0 0 0 44 0 0 41 2
463 1001
126 1001
3 0 10 0 0 0 0 43 0 0 41 2
463 1042
126 1042
3 0 10 0 0 0 0 52 0 0 41 2
461 1349
126 1349
3 0 10 0 0 0 0 55 0 0 41 2
462 1227
126 1227
3 0 10 0 0 0 0 56 0 0 41 2
462 1187
126 1187
4 0 11 0 0 0 0 51 0 0 204 2
461 1399
183 1399
3 0 10 0 0 0 0 51 0 0 41 2
461 1390
126 1390
2 0 10 0 0 4224 0 68 0 0 0 2
126 49
126 1426
4 0 12 0 0 4096 0 52 0 0 211 2
461 1358
146 1358
4 0 11 0 0 0 0 53 0 0 204 2
461 1317
183 1317
3 0 13 0 0 4096 0 53 0 0 210 2
461 1308
91 1308
4 0 12 0 0 0 0 54 0 0 211 2
461 1277
146 1277
3 0 13 0 0 0 0 54 0 0 210 2
461 1268
91 1268
2 0 14 0 0 4096 0 51 0 0 205 2
461 1381
60 1381
2 0 14 0 0 0 0 52 0 0 205 2
461 1340
60 1340
4 0 11 0 0 0 0 55 0 0 204 2
462 1236
183 1236
4 0 12 0 0 4096 0 56 0 0 211 2
462 1196
146 1196
4 0 11 0 0 0 0 57 0 0 204 2
463 1156
183 1156
3 0 13 0 0 4096 0 57 0 0 210 2
463 1147
91 1147
4 0 12 0 0 4096 0 58 0 0 211 2
464 1115
146 1115
3 0 13 0 0 4096 0 58 0 0 210 2
464 1106
91 1106
2 0 14 0 0 0 0 53 0 0 205 2
461 1299
60 1299
2 0 14 0 0 0 0 54 0 0 205 2
461 1259
60 1259
2 0 15 0 0 4096 0 55 0 0 209 2
462 1218
25 1218
2 0 15 0 0 0 0 56 0 0 209 2
462 1178
25 1178
2 0 15 0 0 4096 0 57 0 0 209 2
463 1138
25 1138
2 0 15 0 0 4096 0 58 0 0 209 2
464 1097
25 1097
1 0 6 0 0 0 0 52 0 0 0 2
461 1331
222 1331
1 0 4 0 0 128 0 53 0 0 0 2
461 1290
223 1290
1 0 4 0 0 128 0 55 0 0 0 2
462 1209
219 1209
1 0 2 0 0 128 0 56 0 0 0 2
462 1169
216 1169
4 0 11 0 0 0 0 43 0 0 204 2
463 1051
183 1051
4 0 12 0 0 0 0 44 0 0 211 2
463 1010
146 1010
4 0 11 0 0 0 0 45 0 0 204 2
463 969
183 969
3 0 13 0 0 0 0 45 0 0 210 2
463 960
91 960
4 0 12 0 0 0 0 46 0 0 211 2
463 929
146 929
3 0 13 0 0 0 0 46 0 0 210 2
463 920
91 920
4 0 11 0 0 0 0 47 0 0 204 2
464 888
183 888
4 0 12 0 0 0 0 48 0 0 211 2
464 848
146 848
4 0 11 0 0 0 0 49 0 0 204 2
465 808
183 808
3 0 13 0 0 4096 0 49 0 0 210 2
465 799
91 799
4 0 12 0 0 4096 0 50 0 0 211 2
466 767
146 767
3 0 13 0 0 4096 0 50 0 0 210 2
466 758
91 758
2 0 14 0 0 4096 0 43 0 0 205 2
463 1033
60 1033
2 0 14 0 0 0 0 44 0 0 205 2
463 992
60 992
2 0 14 0 0 0 0 45 0 0 205 2
463 951
60 951
2 0 14 0 0 0 0 46 0 0 205 2
463 911
60 911
2 0 15 0 0 0 0 47 0 0 209 2
464 870
25 870
2 0 15 0 0 0 0 48 0 0 209 2
464 830
25 830
1 0 7 0 0 0 0 44 0 0 0 2
463 983
214 983
1 0 5 0 0 0 0 45 0 0 0 2
463 942
216 942
1 0 3 0 0 128 0 46 0 0 0 2
463 902
217 902
1 0 5 0 0 128 0 47 0 0 0 2
464 861
213 861
1 0 3 0 0 128 0 48 0 0 0 2
464 821
215 821
2 0 15 0 0 4096 0 49 0 0 209 2
465 790
25 790
2 0 15 0 0 4096 0 50 0 0 209 2
466 749
25 749
4 0 12 0 0 0 0 36 0 0 211 2
466 667
146 667
4 0 11 0 0 0 0 37 0 0 204 2
466 626
183 626
3 0 13 0 0 0 0 37 0 0 210 2
466 617
91 617
4 0 12 0 0 0 0 38 0 0 211 2
466 586
146 586
3 0 13 0 0 0 0 38 0 0 210 2
466 577
91 577
2 0 14 0 0 4096 0 35 0 0 205 2
466 690
60 690
2 0 14 0 0 0 0 36 0 0 205 2
466 649
60 649
2 0 14 0 0 0 0 37 0 0 205 2
466 608
60 608
2 0 14 0 0 0 0 38 0 0 205 2
466 568
60 568
1 0 8 0 0 0 0 36 0 0 0 2
466 640
223 640
1 0 2 0 0 0 0 37 0 0 0 2
466 599
219 599
1 0 4 0 0 128 0 38 0 0 0 2
466 559
219 559
4 0 11 0 0 4096 0 39 0 0 204 2
467 545
183 545
2 0 15 0 0 4096 0 39 0 0 209 2
467 527
25 527
1 0 2 0 0 128 0 39 0 0 0 2
467 518
217 518
4 0 12 0 0 4096 0 40 0 0 211 2
467 505
146 505
2 0 15 0 0 0 0 40 0 0 209 2
467 487
25 487
1 0 4 0 0 128 0 40 0 0 0 2
467 478
218 478
0 0 11 0 0 4096 0 0 0 0 204 2
475 465
183 465
3 0 13 0 0 4096 0 41 0 0 210 2
468 456
91 456
2 0 15 0 0 4096 0 41 0 0 209 2
468 447
25 447
4 0 12 0 0 4096 0 42 0 0 211 2
469 424
146 424
3 0 13 0 0 4096 0 42 0 0 210 2
469 415
91 415
2 0 15 0 0 4096 0 42 0 0 209 2
469 406
25 406
4 0 11 0 0 0 0 59 0 0 204 2
469 373
183 373
2 0 14 0 0 4096 0 59 0 0 205 2
469 355
60 355
4 0 12 0 0 0 0 60 0 0 211 2
469 332
146 332
2 0 14 0 0 0 0 60 0 0 205 2
469 314
60 314
1 0 9 0 0 0 0 60 0 0 0 2
469 305
213 305
4 0 11 0 0 0 0 61 0 0 204 2
469 291
183 291
3 0 13 0 0 0 0 61 0 0 210 2
469 282
91 282
2 0 14 0 0 0 0 61 0 0 205 2
469 273
60 273
4 0 12 0 0 0 0 62 0 0 211 2
469 251
146 251
3 0 13 0 0 0 0 62 0 0 210 2
469 242
91 242
2 0 14 0 0 0 0 62 0 0 205 2
469 233
60 233
1 0 5 0 0 128 0 62 0 0 0 2
469 224
212 224
1 0 3 0 0 128 0 63 0 0 0 2
470 183
211 183
1 0 5 0 0 128 0 64 0 0 0 2
470 143
217 143
4 0 15 0 0 4096 0 63 0 0 209 2
470 210
25 210
3 0 11 0 0 0 0 63 0 0 204 2
470 201
183 201
4 0 12 0 0 4096 0 64 0 0 211 2
470 170
146 170
2 0 15 0 0 0 0 64 0 0 209 2
470 152
25 152
4 0 11 0 0 0 0 65 0 0 204 2
471 130
183 130
3 0 13 0 0 4096 0 65 0 0 210 2
471 121
91 121
2 0 15 0 0 4096 0 65 0 0 209 2
471 112
25 112
4 0 12 0 0 4096 0 66 0 0 211 2
472 89
146 89
3 0 13 0 0 4096 0 66 0 0 210 2
472 80
91 80
2 0 15 0 0 4096 0 66 0 0 209 2
472 71
25 71
1 0 16 0 0 4096 0 66 0 0 141 2
472 62
408 62
1 0 16 0 0 0 0 42 0 0 141 2
469 397
408 397
0 1 16 0 0 0 0 0 50 141 0 2
408 740
466 740
1 1 16 0 0 4224 0 2 58 0 0 3
408 47
408 1088
464 1088
1 0 17 0 0 4096 0 57 0 0 146 2
463 1129
375 1129
1 0 17 0 0 4096 0 49 0 0 146 2
465 781
375 781
1 0 17 0 0 4096 0 41 0 0 146 2
468 438
375 438
1 0 17 0 0 4096 0 65 0 0 147 2
471 103
375 103
0 1 17 0 0 4224 0 0 54 147 0 3
375 263
375 1250
461 1250
1 1 17 0 0 0 0 3 61 0 0 3
375 46
375 264
469 264
5 4 18 0 0 4224 0 59 33 0 0 4
514 359
640 359
640 304
644 304
5 3 19 0 0 4224 0 60 33 0 0 4
514 318
629 318
629 295
644 295
5 2 20 0 0 4224 0 61 33 0 0 4
514 277
608 277
608 286
644 286
5 1 21 0 0 4224 0 62 33 0 0 4
514 237
618 237
618 277
644 277
5 4 22 0 0 4224 0 63 34 0 0 3
515 196
657 196
657 133
5 3 23 0 0 4224 0 64 34 0 0 4
515 156
652 156
652 124
657 124
5 2 24 0 0 8320 0 65 34 0 0 3
516 116
516 115
657 115
5 1 25 0 0 8320 0 66 34 0 0 3
517 75
517 106
657 106
5 4 26 0 0 4224 0 39 32 0 0 3
512 531
648 531
648 471
5 3 27 0 0 4224 0 40 32 0 0 4
512 491
628 491
628 462
648 462
5 2 28 0 0 4224 0 41 32 0 0 4
513 451
617 451
617 453
648 453
5 1 29 0 0 4224 0 42 32 0 0 4
514 410
629 410
629 444
648 444
5 1 30 0 0 4224 0 38 15 0 0 4
511 572
631 572
631 609
643 609
5 2 31 0 0 4224 0 37 15 0 0 4
511 612
631 612
631 618
643 618
5 3 32 0 0 4224 0 36 15 0 0 4
511 653
629 653
629 627
643 627
5 4 33 0 0 4224 0 35 15 0 0 3
511 694
643 694
643 636
5 1 34 0 0 4224 0 46 30 0 0 4
508 915
628 915
628 948
650 948
5 4 35 0 0 4224 0 47 31 0 0 4
509 874
629 874
629 818
649 818
5 2 36 0 0 4224 0 45 30 0 0 4
508 955
618 955
618 957
650 957
5 3 37 0 0 4224 0 48 31 0 0 4
509 834
618 834
618 809
649 809
5 3 38 0 0 4224 0 44 30 0 0 4
508 996
617 996
617 966
650 966
5 2 39 0 0 4224 0 49 31 0 0 4
510 794
618 794
618 800
649 800
5 4 40 0 0 4224 0 43 30 0 0 4
508 1037
628 1037
628 975
650 975
5 1 41 0 0 4224 0 50 31 0 0 4
511 753
629 753
629 791
649 791
5 1 42 0 0 4224 0 58 29 0 0 4
509 1101
632 1101
632 1127
652 1127
5 2 43 0 0 4224 0 57 29 0 0 4
508 1142
616 1142
616 1136
652 1136
5 3 44 0 0 4224 0 56 29 0 0 4
507 1182
640 1182
640 1145
652 1145
5 4 45 0 0 4224 0 55 29 0 0 3
507 1222
652 1222
652 1154
5 2 46 0 0 4224 0 53 28 0 0 4
506 1303
612 1303
612 1296
652 1296
5 1 47 0 0 4224 0 54 28 0 0 4
506 1263
621 1263
621 1287
652 1287
5 3 48 0 0 4224 0 52 28 0 0 4
506 1344
619 1344
619 1305
652 1305
5 4 49 0 0 4224 0 51 28 0 0 4
506 1385
632 1385
632 1314
652 1314
2 5 50 0 0 8320 0 20 28 0 0 3
789 1183
702 1183
702 1300
5 1 51 0 0 8320 0 29 20 0 0 3
702 1140
702 1165
789 1165
5 2 52 0 0 8320 0 30 21 0 0 3
700 961
700 879
783 879
5 1 53 0 0 8320 0 31 21 0 0 3
699 804
699 861
783 861
5 2 54 0 0 4224 0 15 22 0 0 3
693 622
693 529
776 529
5 1 55 0 0 8320 0 32 22 0 0 3
698 457
698 511
776 511
5 2 56 0 0 4224 0 33 23 0 0 3
694 290
694 195
775 195
5 1 57 0 0 8320 0 34 23 0 0 3
707 119
707 177
775 177
3 1 58 0 0 12416 0 23 24 0 0 4
821 186
851 186
851 180
952 180
3 1 59 0 0 12416 0 22 25 0 0 4
822 520
837 520
837 507
969 507
3 1 60 0 0 12416 0 21 26 0 0 4
829 870
880 870
880 845
961 845
3 1 61 0 0 4224 0 20 27 0 0 4
835 1174
976 1174
976 1183
984 1183
2 0 62 0 0 4096 0 26 0 0 199 2
961 863
907 863
2 0 62 0 0 4096 0 25 0 0 199 2
969 525
907 525
2 0 62 0 0 0 0 24 0 0 199 2
952 198
907 198
1 3 63 0 0 4224 0 19 27 0 0 3
1227 191
1227 1192
1029 1192
1 3 64 0 0 4224 0 17 25 0 0 3
1142 194
1142 516
1014 516
3 1 65 0 0 8320 0 26 18 0 0 3
1006 854
1189 854
1189 193
3 1 66 0 0 4224 0 24 16 0 0 3
997 189
1107 189
1107 193
1 2 62 0 0 4224 0 1 27 0 0 3
907 45
907 1201
984 1201
1 1 3 0 0 4224 0 4 51 0 0 3
337 47
337 1372
461 1372
1 1 4 0 0 4224 0 5 43 0 0 3
302 47
302 1024
463 1024
1 1 5 0 0 4224 0 6 35 0 0 3
266 47
266 681
466 681
1 1 2 0 0 128 0 59 7 0 0 3
469 346
232 346
232 46
2 0 11 0 0 4224 0 69 0 0 0 2
183 51
183 1452
2 0 14 0 0 4224 0 67 0 0 0 2
60 48
60 1401
1 0 15 0 0 0 0 67 0 0 209 2
24 48
25 48
1 0 13 0 0 0 0 68 0 0 210 2
90 49
91 49
1 0 12 0 0 0 0 69 0 0 211 2
147 51
146 51
1 0 15 0 0 4224 0 8 0 0 0 2
25 47
25 1401
1 0 13 0 0 4224 0 9 0 0 0 2
91 47
91 1402
1 0 12 0 0 4224 0 10 0 0 0 2
146 46
146 1399
32
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
473 1379 492 1395
473 1379 492 1395
2 i0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
477 1031 496 1047
477 1031 496 1047
2 i0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
479 687 498 703
479 687 498 703
2 i0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
484 353 503 369
484 353 503 369
2 i0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
473 1338 492 1354
473 1338 492 1354
2 i1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
475 985 494 1001
475 985 494 1001
2 i1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
481 646 500 662
481 646 500 662
2 i1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
483 309 502 325
483 309 502 325
2 i1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
472 1296 491 1312
472 1296 491 1312
2 i2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
478 947 497 963
478 947 497 963
2 i2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
478 604 497 620
478 604 497 620
2 i2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
479 268 498 284
479 268 498 284
2 i2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
472 1255 491 1271
472 1255 491 1271
2 i3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
478 907 497 923
478 907 497 923
2 i3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
479 563 498 579
479 563 498 579
2 i3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
482 229 501 245
482 229 501 245
2 i3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
473 1214 492 1230
473 1214 492 1230
2 i4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
473 867 492 883
473 867 492 883
2 i4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
480 522 499 538
480 522 499 538
2 i4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
483 188 502 204
483 188 502 204
2 i4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
472 1176 491 1192
472 1176 491 1192
2 i5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
477 825 496 841
477 825 496 841
2 i5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
477 483 496 499
477 483 496 499
2 i5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
482 147 501 163
482 147 501 163
2 i5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
475 1133 494 1149
475 1133 494 1149
2 i6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
477 787 496 803
477 787 496 803
2 i6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
478 442 497 458
478 442 497 458
2 i6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
484 108 503 124
484 108 503 124
2 i6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
476 1094 495 1110
476 1094 495 1110
2 i7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
477 744 496 760
477 744 496 760
2 i7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
482 399 501 415
482 399 501 415
2 i7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
483 66 502 82
483 66 502 82
2 i7
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
